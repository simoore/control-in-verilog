module example_hann_function #
(
    parameter IW = 11,
    parameter OW = 13,
    parameter N_RAM = 1250
)(
    input logic clk,
    input logic ce_in,
    input logic [IW-1:0] sig_in,
    output logic ce_out,
    output logic [OW-1:0] sig_out
);

    logic ce_buf;
    logic [IW-1:0] sig_in_buf;
    logic [OW-1:0] func_lut [0:N_RAM-1];
      
    // Input buffer.
    always_ff @(posedge clk) begin
        ce_buf <= ce_in;
        if(ce_in) sig_in_buf <= sig_in;
    end
    
    // Lookup table read.
    always_ff @(posedge clk) begin
        ce_out <= ce_buf;
        sig_out <= func_lut[sig_in_buf];
    end

    initial begin
        ce_buf = 0;
        sig_in_buf = 0;
         
        func_lut[0] = 3225;  
        func_lut[1] = 3226;  
        func_lut[2] = 3228;  
        func_lut[3] = 3229;  
        func_lut[4] = 3230;  
        func_lut[5] = 3232;  
        func_lut[6] = 3233;  
        func_lut[7] = 3234;  
        func_lut[8] = 3235;  
        func_lut[9] = 3237;  
        func_lut[10] = 3238;  
        func_lut[11] = 3239;  
        func_lut[12] = 3241;  
        func_lut[13] = 3242;  
        func_lut[14] = 3243;  
        func_lut[15] = 3244;  
        func_lut[16] = 3246;  
        func_lut[17] = 3247;  
        func_lut[18] = 3248;  
        func_lut[19] = 3249;  
        func_lut[20] = 3251;  
        func_lut[21] = 3252;  
        func_lut[22] = 3253;  
        func_lut[23] = 3255;  
        func_lut[24] = 3256;  
        func_lut[25] = 3257;  
        func_lut[26] = 3258;  
        func_lut[27] = 3260;  
        func_lut[28] = 3261;  
        func_lut[29] = 3262;  
        func_lut[30] = 3263;  
        func_lut[31] = 3265;  
        func_lut[32] = 3266;  
        func_lut[33] = 3267;  
        func_lut[34] = 3268;  
        func_lut[35] = 3270;  
        func_lut[36] = 3271;  
        func_lut[37] = 3272;  
        func_lut[38] = 3273;  
        func_lut[39] = 3275;  
        func_lut[40] = 3276;  
        func_lut[41] = 3277;  
        func_lut[42] = 3279;  
        func_lut[43] = 3280;  
        func_lut[44] = 3281;  
        func_lut[45] = 3282;  
        func_lut[46] = 3284;  
        func_lut[47] = 3285;  
        func_lut[48] = 3286;  
        func_lut[49] = 3287;  
        func_lut[50] = 3289;  
        func_lut[51] = 3290;  
        func_lut[52] = 3291;  
        func_lut[53] = 3292;  
        func_lut[54] = 3294;  
        func_lut[55] = 3295;  
        func_lut[56] = 3296;  
        func_lut[57] = 3297;  
        func_lut[58] = 3299;  
        func_lut[59] = 3300;  
        func_lut[60] = 3301;  
        func_lut[61] = 3302;  
        func_lut[62] = 3303;  
        func_lut[63] = 3305;  
        func_lut[64] = 3306;  
        func_lut[65] = 3307;  
        func_lut[66] = 3308;  
        func_lut[67] = 3310;  
        func_lut[68] = 3311;  
        func_lut[69] = 3312;  
        func_lut[70] = 3313;  
        func_lut[71] = 3315;  
        func_lut[72] = 3316;  
        func_lut[73] = 3317;  
        func_lut[74] = 3318;  
        func_lut[75] = 3320;  
        func_lut[76] = 3321;  
        func_lut[77] = 3322;  
        func_lut[78] = 3323;  
        func_lut[79] = 3324;  
        func_lut[80] = 3326;  
        func_lut[81] = 3327;  
        func_lut[82] = 3328;  
        func_lut[83] = 3329;  
        func_lut[84] = 3331;  
        func_lut[85] = 3332;  
        func_lut[86] = 3333;  
        func_lut[87] = 3334;  
        func_lut[88] = 3335;  
        func_lut[89] = 3337;  
        func_lut[90] = 3338;  
        func_lut[91] = 3339;  
        func_lut[92] = 3340;  
        func_lut[93] = 3342;  
        func_lut[94] = 3343;  
        func_lut[95] = 3344;  
        func_lut[96] = 3345;  
        func_lut[97] = 3346;  
        func_lut[98] = 3348;  
        func_lut[99] = 3349;  
        func_lut[100] = 3350;  
        func_lut[101] = 3351;  
        func_lut[102] = 3353;  
        func_lut[103] = 3354;  
        func_lut[104] = 3355;  
        func_lut[105] = 3356;  
        func_lut[106] = 3357;  
        func_lut[107] = 3359;  
        func_lut[108] = 3360;  
        func_lut[109] = 3361;  
        func_lut[110] = 3362;  
        func_lut[111] = 3363;  
        func_lut[112] = 3365;  
        func_lut[113] = 3366;  
        func_lut[114] = 3367;  
        func_lut[115] = 3368;  
        func_lut[116] = 3369;  
        func_lut[117] = 3371;  
        func_lut[118] = 3372;  
        func_lut[119] = 3373;  
        func_lut[120] = 3374;  
        func_lut[121] = 3375;  
        func_lut[122] = 3377;  
        func_lut[123] = 3378;  
        func_lut[124] = 3379;  
        func_lut[125] = 3380;  
        func_lut[126] = 3381;  
        func_lut[127] = 3383;  
        func_lut[128] = 3384;  
        func_lut[129] = 3385;  
        func_lut[130] = 3386;  
        func_lut[131] = 3387;  
        func_lut[132] = 3389;  
        func_lut[133] = 3390;  
        func_lut[134] = 3391;  
        func_lut[135] = 3392;  
        func_lut[136] = 3393;  
        func_lut[137] = 3394;  
        func_lut[138] = 3396;  
        func_lut[139] = 3397;  
        func_lut[140] = 3398;  
        func_lut[141] = 3399;  
        func_lut[142] = 3400;  
        func_lut[143] = 3402;  
        func_lut[144] = 3403;  
        func_lut[145] = 3404;  
        func_lut[146] = 3405;  
        func_lut[147] = 3406;  
        func_lut[148] = 3407;  
        func_lut[149] = 3409;  
        func_lut[150] = 3410;  
        func_lut[151] = 3411;  
        func_lut[152] = 3412;  
        func_lut[153] = 3413;  
        func_lut[154] = 3414;  
        func_lut[155] = 3416;  
        func_lut[156] = 3417;  
        func_lut[157] = 3418;  
        func_lut[158] = 3419;  
        func_lut[159] = 3420;  
        func_lut[160] = 3421;  
        func_lut[161] = 3423;  
        func_lut[162] = 3424;  
        func_lut[163] = 3425;  
        func_lut[164] = 3426;  
        func_lut[165] = 3427;  
        func_lut[166] = 3428;  
        func_lut[167] = 3430;  
        func_lut[168] = 3431;  
        func_lut[169] = 3432;  
        func_lut[170] = 3433;  
        func_lut[171] = 3434;  
        func_lut[172] = 3435;  
        func_lut[173] = 3437;  
        func_lut[174] = 3438;  
        func_lut[175] = 3439;  
        func_lut[176] = 3440;  
        func_lut[177] = 3441;  
        func_lut[178] = 3442;  
        func_lut[179] = 3443;  
        func_lut[180] = 3445;  
        func_lut[181] = 3446;  
        func_lut[182] = 3447;  
        func_lut[183] = 3448;  
        func_lut[184] = 3449;  
        func_lut[185] = 3450;  
        func_lut[186] = 3451;  
        func_lut[187] = 3453;  
        func_lut[188] = 3454;  
        func_lut[189] = 3455;  
        func_lut[190] = 3456;  
        func_lut[191] = 3457;  
        func_lut[192] = 3458;  
        func_lut[193] = 3459;  
        func_lut[194] = 3461;  
        func_lut[195] = 3462;  
        func_lut[196] = 3463;  
        func_lut[197] = 3464;  
        func_lut[198] = 3465;  
        func_lut[199] = 3466;  
        func_lut[200] = 3467;  
        func_lut[201] = 3469;  
        func_lut[202] = 3470;  
        func_lut[203] = 3471;  
        func_lut[204] = 3472;  
        func_lut[205] = 3473;  
        func_lut[206] = 3474;  
        func_lut[207] = 3475;  
        func_lut[208] = 3476;  
        func_lut[209] = 3478;  
        func_lut[210] = 3479;  
        func_lut[211] = 3480;  
        func_lut[212] = 3481;  
        func_lut[213] = 3482;  
        func_lut[214] = 3483;  
        func_lut[215] = 3484;  
        func_lut[216] = 3485;  
        func_lut[217] = 3487;  
        func_lut[218] = 3488;  
        func_lut[219] = 3489;  
        func_lut[220] = 3490;  
        func_lut[221] = 3491;  
        func_lut[222] = 3492;  
        func_lut[223] = 3493;  
        func_lut[224] = 3494;  
        func_lut[225] = 3495;  
        func_lut[226] = 3497;  
        func_lut[227] = 3498;  
        func_lut[228] = 3499;  
        func_lut[229] = 3500;  
        func_lut[230] = 3501;  
        func_lut[231] = 3502;  
        func_lut[232] = 3503;  
        func_lut[233] = 3504;  
        func_lut[234] = 3505;  
        func_lut[235] = 3507;  
        func_lut[236] = 3508;  
        func_lut[237] = 3509;  
        func_lut[238] = 3510;  
        func_lut[239] = 3511;  
        func_lut[240] = 3512;  
        func_lut[241] = 3513;  
        func_lut[242] = 3514;  
        func_lut[243] = 3515;  
        func_lut[244] = 3516;  
        func_lut[245] = 3518;  
        func_lut[246] = 3519;  
        func_lut[247] = 3520;  
        func_lut[248] = 3521;  
        func_lut[249] = 3522;  
        func_lut[250] = 3523;  
        func_lut[251] = 3524;  
        func_lut[252] = 3525;  
        func_lut[253] = 3526;  
        func_lut[254] = 3527;  
        func_lut[255] = 3528;  
        func_lut[256] = 3530;  
        func_lut[257] = 3531;  
        func_lut[258] = 3532;  
        func_lut[259] = 3533;  
        func_lut[260] = 3534;  
        func_lut[261] = 3535;  
        func_lut[262] = 3536;  
        func_lut[263] = 3537;  
        func_lut[264] = 3538;  
        func_lut[265] = 3539;  
        func_lut[266] = 3540;  
        func_lut[267] = 3541;  
        func_lut[268] = 3542;  
        func_lut[269] = 3544;  
        func_lut[270] = 3545;  
        func_lut[271] = 3546;  
        func_lut[272] = 3547;  
        func_lut[273] = 3548;  
        func_lut[274] = 3549;  
        func_lut[275] = 3550;  
        func_lut[276] = 3551;  
        func_lut[277] = 3552;  
        func_lut[278] = 3553;  
        func_lut[279] = 3554;  
        func_lut[280] = 3555;  
        func_lut[281] = 3556;  
        func_lut[282] = 3557;  
        func_lut[283] = 3558;  
        func_lut[284] = 3560;  
        func_lut[285] = 3561;  
        func_lut[286] = 3562;  
        func_lut[287] = 3563;  
        func_lut[288] = 3564;  
        func_lut[289] = 3565;  
        func_lut[290] = 3566;  
        func_lut[291] = 3567;  
        func_lut[292] = 3568;  
        func_lut[293] = 3569;  
        func_lut[294] = 3570;  
        func_lut[295] = 3571;  
        func_lut[296] = 3572;  
        func_lut[297] = 3573;  
        func_lut[298] = 3574;  
        func_lut[299] = 3575;  
        func_lut[300] = 3576;  
        func_lut[301] = 3577;  
        func_lut[302] = 3578;  
        func_lut[303] = 3580;  
        func_lut[304] = 3581;  
        func_lut[305] = 3582;  
        func_lut[306] = 3583;  
        func_lut[307] = 3584;  
        func_lut[308] = 3585;  
        func_lut[309] = 3586;  
        func_lut[310] = 3587;  
        func_lut[311] = 3588;  
        func_lut[312] = 3589;  
        func_lut[313] = 3590;  
        func_lut[314] = 3591;  
        func_lut[315] = 3592;  
        func_lut[316] = 3593;  
        func_lut[317] = 3594;  
        func_lut[318] = 3595;  
        func_lut[319] = 3596;  
        func_lut[320] = 3597;  
        func_lut[321] = 3598;  
        func_lut[322] = 3599;  
        func_lut[323] = 3600;  
        func_lut[324] = 3601;  
        func_lut[325] = 3602;  
        func_lut[326] = 3603;  
        func_lut[327] = 3604;  
        func_lut[328] = 3605;  
        func_lut[329] = 3606;  
        func_lut[330] = 3607;  
        func_lut[331] = 3608;  
        func_lut[332] = 3609;  
        func_lut[333] = 3610;  
        func_lut[334] = 3611;  
        func_lut[335] = 3612;  
        func_lut[336] = 3613;  
        func_lut[337] = 3614;  
        func_lut[338] = 3615;  
        func_lut[339] = 3616;  
        func_lut[340] = 3617;  
        func_lut[341] = 3618;  
        func_lut[342] = 3619;  
        func_lut[343] = 3620;  
        func_lut[344] = 3622;  
        func_lut[345] = 3623;  
        func_lut[346] = 3624;  
        func_lut[347] = 3625;  
        func_lut[348] = 3626;  
        func_lut[349] = 3627;  
        func_lut[350] = 3628;  
        func_lut[351] = 3629;  
        func_lut[352] = 3630;  
        func_lut[353] = 3631;  
        func_lut[354] = 3632;  
        func_lut[355] = 3633;  
        func_lut[356] = 3634;  
        func_lut[357] = 3634;  
        func_lut[358] = 3635;  
        func_lut[359] = 3636;  
        func_lut[360] = 3637;  
        func_lut[361] = 3638;  
        func_lut[362] = 3639;  
        func_lut[363] = 3640;  
        func_lut[364] = 3641;  
        func_lut[365] = 3642;  
        func_lut[366] = 3643;  
        func_lut[367] = 3644;  
        func_lut[368] = 3645;  
        func_lut[369] = 3646;  
        func_lut[370] = 3647;  
        func_lut[371] = 3648;  
        func_lut[372] = 3649;  
        func_lut[373] = 3650;  
        func_lut[374] = 3651;  
        func_lut[375] = 3652;  
        func_lut[376] = 3653;  
        func_lut[377] = 3654;  
        func_lut[378] = 3655;  
        func_lut[379] = 3656;  
        func_lut[380] = 3657;  
        func_lut[381] = 3658;  
        func_lut[382] = 3659;  
        func_lut[383] = 3660;  
        func_lut[384] = 3661;  
        func_lut[385] = 3662;  
        func_lut[386] = 3663;  
        func_lut[387] = 3664;  
        func_lut[388] = 3665;  
        func_lut[389] = 3666;  
        func_lut[390] = 3667;  
        func_lut[391] = 3668;  
        func_lut[392] = 3669;  
        func_lut[393] = 3670;  
        func_lut[394] = 3671;  
        func_lut[395] = 3672;  
        func_lut[396] = 3673;  
        func_lut[397] = 3673;  
        func_lut[398] = 3674;  
        func_lut[399] = 3675;  
        func_lut[400] = 3676;  
        func_lut[401] = 3677;  
        func_lut[402] = 3678;  
        func_lut[403] = 3679;  
        func_lut[404] = 3680;  
        func_lut[405] = 3681;  
        func_lut[406] = 3682;  
        func_lut[407] = 3683;  
        func_lut[408] = 3684;  
        func_lut[409] = 3685;  
        func_lut[410] = 3686;  
        func_lut[411] = 3687;  
        func_lut[412] = 3688;  
        func_lut[413] = 3689;  
        func_lut[414] = 3690;  
        func_lut[415] = 3691;  
        func_lut[416] = 3691;  
        func_lut[417] = 3692;  
        func_lut[418] = 3693;  
        func_lut[419] = 3694;  
        func_lut[420] = 3695;  
        func_lut[421] = 3696;  
        func_lut[422] = 3697;  
        func_lut[423] = 3698;  
        func_lut[424] = 3699;  
        func_lut[425] = 3700;  
        func_lut[426] = 3701;  
        func_lut[427] = 3702;  
        func_lut[428] = 3703;  
        func_lut[429] = 3704;  
        func_lut[430] = 3704;  
        func_lut[431] = 3705;  
        func_lut[432] = 3706;  
        func_lut[433] = 3707;  
        func_lut[434] = 3708;  
        func_lut[435] = 3709;  
        func_lut[436] = 3710;  
        func_lut[437] = 3711;  
        func_lut[438] = 3712;  
        func_lut[439] = 3713;  
        func_lut[440] = 3714;  
        func_lut[441] = 3715;  
        func_lut[442] = 3716;  
        func_lut[443] = 3716;  
        func_lut[444] = 3717;  
        func_lut[445] = 3718;  
        func_lut[446] = 3719;  
        func_lut[447] = 3720;  
        func_lut[448] = 3721;  
        func_lut[449] = 3722;  
        func_lut[450] = 3723;  
        func_lut[451] = 3724;  
        func_lut[452] = 3725;  
        func_lut[453] = 3725;  
        func_lut[454] = 3726;  
        func_lut[455] = 3727;  
        func_lut[456] = 3728;  
        func_lut[457] = 3729;  
        func_lut[458] = 3730;  
        func_lut[459] = 3731;  
        func_lut[460] = 3732;  
        func_lut[461] = 3733;  
        func_lut[462] = 3734;  
        func_lut[463] = 3734;  
        func_lut[464] = 3735;  
        func_lut[465] = 3736;  
        func_lut[466] = 3737;  
        func_lut[467] = 3738;  
        func_lut[468] = 3739;  
        func_lut[469] = 3740;  
        func_lut[470] = 3741;  
        func_lut[471] = 3742;  
        func_lut[472] = 3742;  
        func_lut[473] = 3743;  
        func_lut[474] = 3744;  
        func_lut[475] = 3745;  
        func_lut[476] = 3746;  
        func_lut[477] = 3747;  
        func_lut[478] = 3748;  
        func_lut[479] = 3749;  
        func_lut[480] = 3749;  
        func_lut[481] = 3750;  
        func_lut[482] = 3751;  
        func_lut[483] = 3752;  
        func_lut[484] = 3753;  
        func_lut[485] = 3754;  
        func_lut[486] = 3755;  
        func_lut[487] = 3756;  
        func_lut[488] = 3756;  
        func_lut[489] = 3757;  
        func_lut[490] = 3758;  
        func_lut[491] = 3759;  
        func_lut[492] = 3760;  
        func_lut[493] = 3761;  
        func_lut[494] = 3762;  
        func_lut[495] = 3762;  
        func_lut[496] = 3763;  
        func_lut[497] = 3764;  
        func_lut[498] = 3765;  
        func_lut[499] = 3766;  
        func_lut[500] = 3767;  
        func_lut[501] = 3768;  
        func_lut[502] = 3768;  
        func_lut[503] = 3769;  
        func_lut[504] = 3770;  
        func_lut[505] = 3771;  
        func_lut[506] = 3772;  
        func_lut[507] = 3773;  
        func_lut[508] = 3774;  
        func_lut[509] = 3774;  
        func_lut[510] = 3775;  
        func_lut[511] = 3776;  
        func_lut[512] = 3777;  
        func_lut[513] = 3778;  
        func_lut[514] = 3779;  
        func_lut[515] = 3779;  
        func_lut[516] = 3780;  
        func_lut[517] = 3781;  
        func_lut[518] = 3782;  
        func_lut[519] = 3783;  
        func_lut[520] = 3784;  
        func_lut[521] = 3784;  
        func_lut[522] = 3785;  
        func_lut[523] = 3786;  
        func_lut[524] = 3787;  
        func_lut[525] = 3788;  
        func_lut[526] = 3789;  
        func_lut[527] = 3789;  
        func_lut[528] = 3790;  
        func_lut[529] = 3791;  
        func_lut[530] = 3792;  
        func_lut[531] = 3793;  
        func_lut[532] = 3794;  
        func_lut[533] = 3794;  
        func_lut[534] = 3795;  
        func_lut[535] = 3796;  
        func_lut[536] = 3797;  
        func_lut[537] = 3798;  
        func_lut[538] = 3798;  
        func_lut[539] = 3799;  
        func_lut[540] = 3800;  
        func_lut[541] = 3801;  
        func_lut[542] = 3802;  
        func_lut[543] = 3803;  
        func_lut[544] = 3803;  
        func_lut[545] = 3804;  
        func_lut[546] = 3805;  
        func_lut[547] = 3806;  
        func_lut[548] = 3807;  
        func_lut[549] = 3807;  
        func_lut[550] = 3808;  
        func_lut[551] = 3809;  
        func_lut[552] = 3810;  
        func_lut[553] = 3811;  
        func_lut[554] = 3811;  
        func_lut[555] = 3812;  
        func_lut[556] = 3813;  
        func_lut[557] = 3814;  
        func_lut[558] = 3815;  
        func_lut[559] = 3815;  
        func_lut[560] = 3816;  
        func_lut[561] = 3817;  
        func_lut[562] = 3818;  
        func_lut[563] = 3819;  
        func_lut[564] = 3819;  
        func_lut[565] = 3820;  
        func_lut[566] = 3821;  
        func_lut[567] = 3822;  
        func_lut[568] = 3822;  
        func_lut[569] = 3823;  
        func_lut[570] = 3824;  
        func_lut[571] = 3825;  
        func_lut[572] = 3826;  
        func_lut[573] = 3826;  
        func_lut[574] = 3827;  
        func_lut[575] = 3828;  
        func_lut[576] = 3829;  
        func_lut[577] = 3829;  
        func_lut[578] = 3830;  
        func_lut[579] = 3831;  
        func_lut[580] = 3832;  
        func_lut[581] = 3833;  
        func_lut[582] = 3833;  
        func_lut[583] = 3834;  
        func_lut[584] = 3835;  
        func_lut[585] = 3836;  
        func_lut[586] = 3836;  
        func_lut[587] = 3837;  
        func_lut[588] = 3838;  
        func_lut[589] = 3839;  
        func_lut[590] = 3839;  
        func_lut[591] = 3840;  
        func_lut[592] = 3841;  
        func_lut[593] = 3842;  
        func_lut[594] = 3843;  
        func_lut[595] = 3843;  
        func_lut[596] = 3844;  
        func_lut[597] = 3845;  
        func_lut[598] = 3846;  
        func_lut[599] = 3846;  
        func_lut[600] = 3847;  
        func_lut[601] = 3848;  
        func_lut[602] = 3849;  
        func_lut[603] = 3849;  
        func_lut[604] = 3850;  
        func_lut[605] = 3851;  
        func_lut[606] = 3852;  
        func_lut[607] = 3852;  
        func_lut[608] = 3853;  
        func_lut[609] = 3854;  
        func_lut[610] = 3854;  
        func_lut[611] = 3855;  
        func_lut[612] = 3856;  
        func_lut[613] = 3857;  
        func_lut[614] = 3857;  
        func_lut[615] = 3858;  
        func_lut[616] = 3859;  
        func_lut[617] = 3860;  
        func_lut[618] = 3860;  
        func_lut[619] = 3861;  
        func_lut[620] = 3862;  
        func_lut[621] = 3863;  
        func_lut[622] = 3863;  
        func_lut[623] = 3864;  
        func_lut[624] = 3865;  
        func_lut[625] = 3865;  
        func_lut[626] = 3866;  
        func_lut[627] = 3867;  
        func_lut[628] = 3868;  
        func_lut[629] = 3868;  
        func_lut[630] = 3869;  
        func_lut[631] = 3870;  
        func_lut[632] = 3871;  
        func_lut[633] = 3871;  
        func_lut[634] = 3872;  
        func_lut[635] = 3873;  
        func_lut[636] = 3873;  
        func_lut[637] = 3874;  
        func_lut[638] = 3875;  
        func_lut[639] = 3876;  
        func_lut[640] = 3876;  
        func_lut[641] = 3877;  
        func_lut[642] = 3878;  
        func_lut[643] = 3878;  
        func_lut[644] = 3879;  
        func_lut[645] = 3880;  
        func_lut[646] = 3880;  
        func_lut[647] = 3881;  
        func_lut[648] = 3882;  
        func_lut[649] = 3883;  
        func_lut[650] = 3883;  
        func_lut[651] = 3884;  
        func_lut[652] = 3885;  
        func_lut[653] = 3885;  
        func_lut[654] = 3886;  
        func_lut[655] = 3887;  
        func_lut[656] = 3887;  
        func_lut[657] = 3888;  
        func_lut[658] = 3889;  
        func_lut[659] = 3889;  
        func_lut[660] = 3890;  
        func_lut[661] = 3891;  
        func_lut[662] = 3892;  
        func_lut[663] = 3892;  
        func_lut[664] = 3893;  
        func_lut[665] = 3894;  
        func_lut[666] = 3894;  
        func_lut[667] = 3895;  
        func_lut[668] = 3896;  
        func_lut[669] = 3896;  
        func_lut[670] = 3897;  
        func_lut[671] = 3898;  
        func_lut[672] = 3898;  
        func_lut[673] = 3899;  
        func_lut[674] = 3900;  
        func_lut[675] = 3900;  
        func_lut[676] = 3901;  
        func_lut[677] = 3902;  
        func_lut[678] = 3902;  
        func_lut[679] = 3903;  
        func_lut[680] = 3904;  
        func_lut[681] = 3904;  
        func_lut[682] = 3905;  
        func_lut[683] = 3906;  
        func_lut[684] = 3906;  
        func_lut[685] = 3907;  
        func_lut[686] = 3908;  
        func_lut[687] = 3908;  
        func_lut[688] = 3909;  
        func_lut[689] = 3910;  
        func_lut[690] = 3910;  
        func_lut[691] = 3911;  
        func_lut[692] = 3912;  
        func_lut[693] = 3912;  
        func_lut[694] = 3913;  
        func_lut[695] = 3914;  
        func_lut[696] = 3914;  
        func_lut[697] = 3915;  
        func_lut[698] = 3915;  
        func_lut[699] = 3916;  
        func_lut[700] = 3917;  
        func_lut[701] = 3917;  
        func_lut[702] = 3918;  
        func_lut[703] = 3919;  
        func_lut[704] = 3919;  
        func_lut[705] = 3920;  
        func_lut[706] = 3921;  
        func_lut[707] = 3921;  
        func_lut[708] = 3922;  
        func_lut[709] = 3922;  
        func_lut[710] = 3923;  
        func_lut[711] = 3924;  
        func_lut[712] = 3924;  
        func_lut[713] = 3925;  
        func_lut[714] = 3926;  
        func_lut[715] = 3926;  
        func_lut[716] = 3927;  
        func_lut[717] = 3928;  
        func_lut[718] = 3928;  
        func_lut[719] = 3929;  
        func_lut[720] = 3929;  
        func_lut[721] = 3930;  
        func_lut[722] = 3931;  
        func_lut[723] = 3931;  
        func_lut[724] = 3932;  
        func_lut[725] = 3932;  
        func_lut[726] = 3933;  
        func_lut[727] = 3934;  
        func_lut[728] = 3934;  
        func_lut[729] = 3935;  
        func_lut[730] = 3936;  
        func_lut[731] = 3936;  
        func_lut[732] = 3937;  
        func_lut[733] = 3937;  
        func_lut[734] = 3938;  
        func_lut[735] = 3939;  
        func_lut[736] = 3939;  
        func_lut[737] = 3940;  
        func_lut[738] = 3940;  
        func_lut[739] = 3941;  
        func_lut[740] = 3942;  
        func_lut[741] = 3942;  
        func_lut[742] = 3943;  
        func_lut[743] = 3943;  
        func_lut[744] = 3944;  
        func_lut[745] = 3945;  
        func_lut[746] = 3945;  
        func_lut[747] = 3946;  
        func_lut[748] = 3946;  
        func_lut[749] = 3947;  
        func_lut[750] = 3947;  
        func_lut[751] = 3948;  
        func_lut[752] = 3949;  
        func_lut[753] = 3949;  
        func_lut[754] = 3950;  
        func_lut[755] = 3950;  
        func_lut[756] = 3951;  
        func_lut[757] = 3952;  
        func_lut[758] = 3952;  
        func_lut[759] = 3953;  
        func_lut[760] = 3953;  
        func_lut[761] = 3954;  
        func_lut[762] = 3954;  
        func_lut[763] = 3955;  
        func_lut[764] = 3956;  
        func_lut[765] = 3956;  
        func_lut[766] = 3957;  
        func_lut[767] = 3957;  
        func_lut[768] = 3958;  
        func_lut[769] = 3958;  
        func_lut[770] = 3959;  
        func_lut[771] = 3960;  
        func_lut[772] = 3960;  
        func_lut[773] = 3961;  
        func_lut[774] = 3961;  
        func_lut[775] = 3962;  
        func_lut[776] = 3962;  
        func_lut[777] = 3963;  
        func_lut[778] = 3964;  
        func_lut[779] = 3964;  
        func_lut[780] = 3965;  
        func_lut[781] = 3965;  
        func_lut[782] = 3966;  
        func_lut[783] = 3966;  
        func_lut[784] = 3967;  
        func_lut[785] = 3967;  
        func_lut[786] = 3968;  
        func_lut[787] = 3968;  
        func_lut[788] = 3969;  
        func_lut[789] = 3970;  
        func_lut[790] = 3970;  
        func_lut[791] = 3971;  
        func_lut[792] = 3971;  
        func_lut[793] = 3972;  
        func_lut[794] = 3972;  
        func_lut[795] = 3973;  
        func_lut[796] = 3973;  
        func_lut[797] = 3974;  
        func_lut[798] = 3974;  
        func_lut[799] = 3975;  
        func_lut[800] = 3975;  
        func_lut[801] = 3976;  
        func_lut[802] = 3977;  
        func_lut[803] = 3977;  
        func_lut[804] = 3978;  
        func_lut[805] = 3978;  
        func_lut[806] = 3979;  
        func_lut[807] = 3979;  
        func_lut[808] = 3980;  
        func_lut[809] = 3980;  
        func_lut[810] = 3981;  
        func_lut[811] = 3981;  
        func_lut[812] = 3982;  
        func_lut[813] = 3982;  
        func_lut[814] = 3983;  
        func_lut[815] = 3983;  
        func_lut[816] = 3984;  
        func_lut[817] = 3984;  
        func_lut[818] = 3985;  
        func_lut[819] = 3985;  
        func_lut[820] = 3986;  
        func_lut[821] = 3986;  
        func_lut[822] = 3987;  
        func_lut[823] = 3987;  
        func_lut[824] = 3988;  
        func_lut[825] = 3988;  
        func_lut[826] = 3989;  
        func_lut[827] = 3989;  
        func_lut[828] = 3990;  
        func_lut[829] = 3990;  
        func_lut[830] = 3991;  
        func_lut[831] = 3991;  
        func_lut[832] = 3992;  
        func_lut[833] = 3992;  
        func_lut[834] = 3993;  
        func_lut[835] = 3993;  
        func_lut[836] = 3994;  
        func_lut[837] = 3994;  
        func_lut[838] = 3995;  
        func_lut[839] = 3995;  
        func_lut[840] = 3996;  
        func_lut[841] = 3996;  
        func_lut[842] = 3997;  
        func_lut[843] = 3997;  
        func_lut[844] = 3998;  
        func_lut[845] = 3998;  
        func_lut[846] = 3999;  
        func_lut[847] = 3999;  
        func_lut[848] = 4000;  
        func_lut[849] = 4000;  
        func_lut[850] = 4001;  
        func_lut[851] = 4001;  
        func_lut[852] = 4002;  
        func_lut[853] = 4002;  
        func_lut[854] = 4002;  
        func_lut[855] = 4003;  
        func_lut[856] = 4003;  
        func_lut[857] = 4004;  
        func_lut[858] = 4004;  
        func_lut[859] = 4005;  
        func_lut[860] = 4005;  
        func_lut[861] = 4006;  
        func_lut[862] = 4006;  
        func_lut[863] = 4007;  
        func_lut[864] = 4007;  
        func_lut[865] = 4008;  
        func_lut[866] = 4008;  
        func_lut[867] = 4008;  
        func_lut[868] = 4009;  
        func_lut[869] = 4009;  
        func_lut[870] = 4010;  
        func_lut[871] = 4010;  
        func_lut[872] = 4011;  
        func_lut[873] = 4011;  
        func_lut[874] = 4012;  
        func_lut[875] = 4012;  
        func_lut[876] = 4013;  
        func_lut[877] = 4013;  
        func_lut[878] = 4013;  
        func_lut[879] = 4014;  
        func_lut[880] = 4014;  
        func_lut[881] = 4015;  
        func_lut[882] = 4015;  
        func_lut[883] = 4016;  
        func_lut[884] = 4016;  
        func_lut[885] = 4016;  
        func_lut[886] = 4017;  
        func_lut[887] = 4017;  
        func_lut[888] = 4018;  
        func_lut[889] = 4018;  
        func_lut[890] = 4019;  
        func_lut[891] = 4019;  
        func_lut[892] = 4019;  
        func_lut[893] = 4020;  
        func_lut[894] = 4020;  
        func_lut[895] = 4021;  
        func_lut[896] = 4021;  
        func_lut[897] = 4022;  
        func_lut[898] = 4022;  
        func_lut[899] = 4022;  
        func_lut[900] = 4023;  
        func_lut[901] = 4023;  
        func_lut[902] = 4024;  
        func_lut[903] = 4024;  
        func_lut[904] = 4024;  
        func_lut[905] = 4025;  
        func_lut[906] = 4025;  
        func_lut[907] = 4026;  
        func_lut[908] = 4026;  
        func_lut[909] = 4027;  
        func_lut[910] = 4027;  
        func_lut[911] = 4027;  
        func_lut[912] = 4028;  
        func_lut[913] = 4028;  
        func_lut[914] = 4029;  
        func_lut[915] = 4029;  
        func_lut[916] = 4029;  
        func_lut[917] = 4030;  
        func_lut[918] = 4030;  
        func_lut[919] = 4031;  
        func_lut[920] = 4031;  
        func_lut[921] = 4031;  
        func_lut[922] = 4032;  
        func_lut[923] = 4032;  
        func_lut[924] = 4032;  
        func_lut[925] = 4033;  
        func_lut[926] = 4033;  
        func_lut[927] = 4034;  
        func_lut[928] = 4034;  
        func_lut[929] = 4034;  
        func_lut[930] = 4035;  
        func_lut[931] = 4035;  
        func_lut[932] = 4036;  
        func_lut[933] = 4036;  
        func_lut[934] = 4036;  
        func_lut[935] = 4037;  
        func_lut[936] = 4037;  
        func_lut[937] = 4037;  
        func_lut[938] = 4038;  
        func_lut[939] = 4038;  
        func_lut[940] = 4039;  
        func_lut[941] = 4039;  
        func_lut[942] = 4039;  
        func_lut[943] = 4040;  
        func_lut[944] = 4040;  
        func_lut[945] = 4040;  
        func_lut[946] = 4041;  
        func_lut[947] = 4041;  
        func_lut[948] = 4041;  
        func_lut[949] = 4042;  
        func_lut[950] = 4042;  
        func_lut[951] = 4043;  
        func_lut[952] = 4043;  
        func_lut[953] = 4043;  
        func_lut[954] = 4044;  
        func_lut[955] = 4044;  
        func_lut[956] = 4044;  
        func_lut[957] = 4045;  
        func_lut[958] = 4045;  
        func_lut[959] = 4045;  
        func_lut[960] = 4046;  
        func_lut[961] = 4046;  
        func_lut[962] = 4046;  
        func_lut[963] = 4047;  
        func_lut[964] = 4047;  
        func_lut[965] = 4047;  
        func_lut[966] = 4048;  
        func_lut[967] = 4048;  
        func_lut[968] = 4048;  
        func_lut[969] = 4049;  
        func_lut[970] = 4049;  
        func_lut[971] = 4049;  
        func_lut[972] = 4050;  
        func_lut[973] = 4050;  
        func_lut[974] = 4050;  
        func_lut[975] = 4051;  
        func_lut[976] = 4051;  
        func_lut[977] = 4051;  
        func_lut[978] = 4052;  
        func_lut[979] = 4052;  
        func_lut[980] = 4052;  
        func_lut[981] = 4053;  
        func_lut[982] = 4053;  
        func_lut[983] = 4053;  
        func_lut[984] = 4054;  
        func_lut[985] = 4054;  
        func_lut[986] = 4054;  
        func_lut[987] = 4055;  
        func_lut[988] = 4055;  
        func_lut[989] = 4055;  
        func_lut[990] = 4056;  
        func_lut[991] = 4056;  
        func_lut[992] = 4056;  
        func_lut[993] = 4056;  
        func_lut[994] = 4057;  
        func_lut[995] = 4057;  
        func_lut[996] = 4057;  
        func_lut[997] = 4058;  
        func_lut[998] = 4058;  
        func_lut[999] = 4058;  
        func_lut[1000] = 4059;  
        func_lut[1001] = 4059;  
        func_lut[1002] = 4059;  
        func_lut[1003] = 4059;  
        func_lut[1004] = 4060;  
        func_lut[1005] = 4060;  
        func_lut[1006] = 4060;  
        func_lut[1007] = 4061;  
        func_lut[1008] = 4061;  
        func_lut[1009] = 4061;  
        func_lut[1010] = 4062;  
        func_lut[1011] = 4062;  
        func_lut[1012] = 4062;  
        func_lut[1013] = 4062;  
        func_lut[1014] = 4063;  
        func_lut[1015] = 4063;  
        func_lut[1016] = 4063;  
        func_lut[1017] = 4064;  
        func_lut[1018] = 4064;  
        func_lut[1019] = 4064;  
        func_lut[1020] = 4064;  
        func_lut[1021] = 4065;  
        func_lut[1022] = 4065;  
        func_lut[1023] = 4065;  
        func_lut[1024] = 4065;  
        func_lut[1025] = 4066;  
        func_lut[1026] = 4066;  
        func_lut[1027] = 4066;  
        func_lut[1028] = 4067;  
        func_lut[1029] = 4067;  
        func_lut[1030] = 4067;  
        func_lut[1031] = 4067;  
        func_lut[1032] = 4068;  
        func_lut[1033] = 4068;  
        func_lut[1034] = 4068;  
        func_lut[1035] = 4068;  
        func_lut[1036] = 4069;  
        func_lut[1037] = 4069;  
        func_lut[1038] = 4069;  
        func_lut[1039] = 4069;  
        func_lut[1040] = 4070;  
        func_lut[1041] = 4070;  
        func_lut[1042] = 4070;  
        func_lut[1043] = 4070;  
        func_lut[1044] = 4071;  
        func_lut[1045] = 4071;  
        func_lut[1046] = 4071;  
        func_lut[1047] = 4071;  
        func_lut[1048] = 4072;  
        func_lut[1049] = 4072;  
        func_lut[1050] = 4072;  
        func_lut[1051] = 4072;  
        func_lut[1052] = 4073;  
        func_lut[1053] = 4073;  
        func_lut[1054] = 4073;  
        func_lut[1055] = 4073;  
        func_lut[1056] = 4073;  
        func_lut[1057] = 4074;  
        func_lut[1058] = 4074;  
        func_lut[1059] = 4074;  
        func_lut[1060] = 4074;  
        func_lut[1061] = 4075;  
        func_lut[1062] = 4075;  
        func_lut[1063] = 4075;  
        func_lut[1064] = 4075;  
        func_lut[1065] = 4076;  
        func_lut[1066] = 4076;  
        func_lut[1067] = 4076;  
        func_lut[1068] = 4076;  
        func_lut[1069] = 4076;  
        func_lut[1070] = 4077;  
        func_lut[1071] = 4077;  
        func_lut[1072] = 4077;  
        func_lut[1073] = 4077;  
        func_lut[1074] = 4077;  
        func_lut[1075] = 4078;  
        func_lut[1076] = 4078;  
        func_lut[1077] = 4078;  
        func_lut[1078] = 4078;  
        func_lut[1079] = 4079;  
        func_lut[1080] = 4079;  
        func_lut[1081] = 4079;  
        func_lut[1082] = 4079;  
        func_lut[1083] = 4079;  
        func_lut[1084] = 4080;  
        func_lut[1085] = 4080;  
        func_lut[1086] = 4080;  
        func_lut[1087] = 4080;  
        func_lut[1088] = 4080;  
        func_lut[1089] = 4080;  
        func_lut[1090] = 4081;  
        func_lut[1091] = 4081;  
        func_lut[1092] = 4081;  
        func_lut[1093] = 4081;  
        func_lut[1094] = 4081;  
        func_lut[1095] = 4082;  
        func_lut[1096] = 4082;  
        func_lut[1097] = 4082;  
        func_lut[1098] = 4082;  
        func_lut[1099] = 4082;  
        func_lut[1100] = 4083;  
        func_lut[1101] = 4083;  
        func_lut[1102] = 4083;  
        func_lut[1103] = 4083;  
        func_lut[1104] = 4083;  
        func_lut[1105] = 4083;  
        func_lut[1106] = 4084;  
        func_lut[1107] = 4084;  
        func_lut[1108] = 4084;  
        func_lut[1109] = 4084;  
        func_lut[1110] = 4084;  
        func_lut[1111] = 4084;  
        func_lut[1112] = 4085;  
        func_lut[1113] = 4085;  
        func_lut[1114] = 4085;  
        func_lut[1115] = 4085;  
        func_lut[1116] = 4085;  
        func_lut[1117] = 4085;  
        func_lut[1118] = 4086;  
        func_lut[1119] = 4086;  
        func_lut[1120] = 4086;  
        func_lut[1121] = 4086;  
        func_lut[1122] = 4086;  
        func_lut[1123] = 4086;  
        func_lut[1124] = 4087;  
        func_lut[1125] = 4087;  
        func_lut[1126] = 4087;  
        func_lut[1127] = 4087;  
        func_lut[1128] = 4087;  
        func_lut[1129] = 4087;  
        func_lut[1130] = 4087;  
        func_lut[1131] = 4088;  
        func_lut[1132] = 4088;  
        func_lut[1133] = 4088;  
        func_lut[1134] = 4088;  
        func_lut[1135] = 4088;  
        func_lut[1136] = 4088;  
        func_lut[1137] = 4088;  
        func_lut[1138] = 4089;  
        func_lut[1139] = 4089;  
        func_lut[1140] = 4089;  
        func_lut[1141] = 4089;  
        func_lut[1142] = 4089;  
        func_lut[1143] = 4089;  
        func_lut[1144] = 4089;  
        func_lut[1145] = 4089;  
        func_lut[1146] = 4090;  
        func_lut[1147] = 4090;  
        func_lut[1148] = 4090;  
        func_lut[1149] = 4090;  
        func_lut[1150] = 4090;  
        func_lut[1151] = 4090;  
        func_lut[1152] = 4090;  
        func_lut[1153] = 4090;  
        func_lut[1154] = 4091;  
        func_lut[1155] = 4091;  
        func_lut[1156] = 4091;  
        func_lut[1157] = 4091;  
        func_lut[1158] = 4091;  
        func_lut[1159] = 4091;  
        func_lut[1160] = 4091;  
        func_lut[1161] = 4091;  
        func_lut[1162] = 4091;  
        func_lut[1163] = 4091;  
        func_lut[1164] = 4092;  
        func_lut[1165] = 4092;  
        func_lut[1166] = 4092;  
        func_lut[1167] = 4092;  
        func_lut[1168] = 4092;  
        func_lut[1169] = 4092;  
        func_lut[1170] = 4092;  
        func_lut[1171] = 4092;  
        func_lut[1172] = 4092;  
        func_lut[1173] = 4092;  
        func_lut[1174] = 4093;  
        func_lut[1175] = 4093;  
        func_lut[1176] = 4093;  
        func_lut[1177] = 4093;  
        func_lut[1178] = 4093;  
        func_lut[1179] = 4093;  
        func_lut[1180] = 4093;  
        func_lut[1181] = 4093;  
        func_lut[1182] = 4093;  
        func_lut[1183] = 4093;  
        func_lut[1184] = 4093;  
        func_lut[1185] = 4093;  
        func_lut[1186] = 4094;  
        func_lut[1187] = 4094;  
        func_lut[1188] = 4094;  
        func_lut[1189] = 4094;  
        func_lut[1190] = 4094;  
        func_lut[1191] = 4094;  
        func_lut[1192] = 4094;  
        func_lut[1193] = 4094;  
        func_lut[1194] = 4094;  
        func_lut[1195] = 4094;  
        func_lut[1196] = 4094;  
        func_lut[1197] = 4094;  
        func_lut[1198] = 4094;  
        func_lut[1199] = 4094;  
        func_lut[1200] = 4095;  
        func_lut[1201] = 4095;  
        func_lut[1202] = 4095;  
        func_lut[1203] = 4095;  
        func_lut[1204] = 4095;  
        func_lut[1205] = 4095;  
        func_lut[1206] = 4095;  
        func_lut[1207] = 4095;  
        func_lut[1208] = 4095;  
        func_lut[1209] = 4095;  
        func_lut[1210] = 4095;  
        func_lut[1211] = 4095;  
        func_lut[1212] = 4095;  
        func_lut[1213] = 4095;  
        func_lut[1214] = 4095;  
        func_lut[1215] = 4095;  
        func_lut[1216] = 4095;  
        func_lut[1217] = 4095;  
        func_lut[1218] = 4095;  
        func_lut[1219] = 4095;  
        func_lut[1220] = 4095;  
        func_lut[1221] = 4096;  
        func_lut[1222] = 4096;  
        func_lut[1223] = 4096;  
        func_lut[1224] = 4096;  
        func_lut[1225] = 4096;  
        func_lut[1226] = 4096;  
        func_lut[1227] = 4096;  
        func_lut[1228] = 4096;  
        func_lut[1229] = 4096;  
        func_lut[1230] = 4096;  
        func_lut[1231] = 4096;  
        func_lut[1232] = 4096;  
        func_lut[1233] = 4096;  
        func_lut[1234] = 4096;  
        func_lut[1235] = 4096;  
        func_lut[1236] = 4096;  
        func_lut[1237] = 4096;  
        func_lut[1238] = 4096;  
        func_lut[1239] = 4096;  
        func_lut[1240] = 4096;  
        func_lut[1241] = 4096;  
        func_lut[1242] = 4096;  
        func_lut[1243] = 4096;  
        func_lut[1244] = 4096;  
        func_lut[1245] = 4096;  
        func_lut[1246] = 4096;  
        func_lut[1247] = 4096;  
        func_lut[1248] = 4096;  
        func_lut[1249] = 4096; 
    end

endmodule