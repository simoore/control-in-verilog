module tree_adder # 
(
)
(
);