module example_nonlinear_function #
(
    parameter IW = 11,
    parameter OW = 14,
    parameter N_RAM = 2048
)(
    input clk,
    input ce_in,
    input [IW-1:0] sig_in,
    output reg ce_out,
    output reg [OW-1:0] sig_out
);

    reg ce_buf;
    reg [IW-1:0] sig_in_buf;
    reg [OW-1:0] func_lut [0:N_RAM-1];
      
    // Input buffer.
    always @(posedge clk) begin
        ce_buf <= ce_in;
        if(ce_in) sig_in_buf <= sig_in;
    end
    
    // Lookup table read.
    always @(posedge clk) begin
        ce_out <= ce_buf;
        sig_out <= func_lut[sig_in_buf];
    end

    initial begin
        ce_buf = 0;
        sig_in_buf = 0;
         
        func_lut[0] = 271;  
        func_lut[1] = 270;  
        func_lut[2] = 270;  
        func_lut[3] = 269;  
        func_lut[4] = 269;  
        func_lut[5] = 269;  
        func_lut[6] = 268;  
        func_lut[7] = 268;  
        func_lut[8] = 267;  
        func_lut[9] = 267;  
        func_lut[10] = 266;  
        func_lut[11] = 266;  
        func_lut[12] = 266;  
        func_lut[13] = 265;  
        func_lut[14] = 265;  
        func_lut[15] = 264;  
        func_lut[16] = 264;  
        func_lut[17] = 264;  
        func_lut[18] = 263;  
        func_lut[19] = 263;  
        func_lut[20] = 262;  
        func_lut[21] = 262;  
        func_lut[22] = 261;  
        func_lut[23] = 261;  
        func_lut[24] = 261;  
        func_lut[25] = 260;  
        func_lut[26] = 260;  
        func_lut[27] = 259;  
        func_lut[28] = 259;  
        func_lut[29] = 259;  
        func_lut[30] = 258;  
        func_lut[31] = 258;  
        func_lut[32] = 257;  
        func_lut[33] = 257;  
        func_lut[34] = 257;  
        func_lut[35] = 256;  
        func_lut[36] = 256;  
        func_lut[37] = 255;  
        func_lut[38] = 255;  
        func_lut[39] = 255;  
        func_lut[40] = 254;  
        func_lut[41] = 254;  
        func_lut[42] = 253;  
        func_lut[43] = 253;  
        func_lut[44] = 253;  
        func_lut[45] = 252;  
        func_lut[46] = 252;  
        func_lut[47] = 251;  
        func_lut[48] = 251;  
        func_lut[49] = 251;  
        func_lut[50] = 250;  
        func_lut[51] = 250;  
        func_lut[52] = 250;  
        func_lut[53] = 249;  
        func_lut[54] = 249;  
        func_lut[55] = 248;  
        func_lut[56] = 248;  
        func_lut[57] = 248;  
        func_lut[58] = 247;  
        func_lut[59] = 247;  
        func_lut[60] = 247;  
        func_lut[61] = 246;  
        func_lut[62] = 246;  
        func_lut[63] = 245;  
        func_lut[64] = 245;  
        func_lut[65] = 245;  
        func_lut[66] = 244;  
        func_lut[67] = 244;  
        func_lut[68] = 244;  
        func_lut[69] = 243;  
        func_lut[70] = 243;  
        func_lut[71] = 242;  
        func_lut[72] = 242;  
        func_lut[73] = 242;  
        func_lut[74] = 241;  
        func_lut[75] = 241;  
        func_lut[76] = 241;  
        func_lut[77] = 240;  
        func_lut[78] = 240;  
        func_lut[79] = 240;  
        func_lut[80] = 239;  
        func_lut[81] = 239;  
        func_lut[82] = 238;  
        func_lut[83] = 238;  
        func_lut[84] = 238;  
        func_lut[85] = 237;  
        func_lut[86] = 237;  
        func_lut[87] = 237;  
        func_lut[88] = 236;  
        func_lut[89] = 236;  
        func_lut[90] = 236;  
        func_lut[91] = 235;  
        func_lut[92] = 235;  
        func_lut[93] = 235;  
        func_lut[94] = 234;  
        func_lut[95] = 234;  
        func_lut[96] = 234;  
        func_lut[97] = 233;  
        func_lut[98] = 233;  
        func_lut[99] = 232;  
        func_lut[100] = 232;  
        func_lut[101] = 232;  
        func_lut[102] = 231;  
        func_lut[103] = 231;  
        func_lut[104] = 231;  
        func_lut[105] = 230;  
        func_lut[106] = 230;  
        func_lut[107] = 230;  
        func_lut[108] = 229;  
        func_lut[109] = 229;  
        func_lut[110] = 229;  
        func_lut[111] = 228;  
        func_lut[112] = 228;  
        func_lut[113] = 228;  
        func_lut[114] = 227;  
        func_lut[115] = 227;  
        func_lut[116] = 227;  
        func_lut[117] = 226;  
        func_lut[118] = 226;  
        func_lut[119] = 226;  
        func_lut[120] = 225;  
        func_lut[121] = 225;  
        func_lut[122] = 225;  
        func_lut[123] = 224;  
        func_lut[124] = 224;  
        func_lut[125] = 224;  
        func_lut[126] = 223;  
        func_lut[127] = 223;  
        func_lut[128] = 223;  
        func_lut[129] = 223;  
        func_lut[130] = 222;  
        func_lut[131] = 222;  
        func_lut[132] = 222;  
        func_lut[133] = 221;  
        func_lut[134] = 221;  
        func_lut[135] = 221;  
        func_lut[136] = 220;  
        func_lut[137] = 220;  
        func_lut[138] = 220;  
        func_lut[139] = 219;  
        func_lut[140] = 219;  
        func_lut[141] = 219;  
        func_lut[142] = 218;  
        func_lut[143] = 218;  
        func_lut[144] = 218;  
        func_lut[145] = 217;  
        func_lut[146] = 217;  
        func_lut[147] = 217;  
        func_lut[148] = 217;  
        func_lut[149] = 216;  
        func_lut[150] = 216;  
        func_lut[151] = 216;  
        func_lut[152] = 215;  
        func_lut[153] = 215;  
        func_lut[154] = 215;  
        func_lut[155] = 214;  
        func_lut[156] = 214;  
        func_lut[157] = 214;  
        func_lut[158] = 213;  
        func_lut[159] = 213;  
        func_lut[160] = 213;  
        func_lut[161] = 213;  
        func_lut[162] = 212;  
        func_lut[163] = 212;  
        func_lut[164] = 212;  
        func_lut[165] = 211;  
        func_lut[166] = 211;  
        func_lut[167] = 211;  
        func_lut[168] = 210;  
        func_lut[169] = 210;  
        func_lut[170] = 210;  
        func_lut[171] = 210;  
        func_lut[172] = 209;  
        func_lut[173] = 209;  
        func_lut[174] = 209;  
        func_lut[175] = 208;  
        func_lut[176] = 208;  
        func_lut[177] = 208;  
        func_lut[178] = 208;  
        func_lut[179] = 207;  
        func_lut[180] = 207;  
        func_lut[181] = 207;  
        func_lut[182] = 206;  
        func_lut[183] = 206;  
        func_lut[184] = 206;  
        func_lut[185] = 205;  
        func_lut[186] = 205;  
        func_lut[187] = 205;  
        func_lut[188] = 205;  
        func_lut[189] = 204;  
        func_lut[190] = 204;  
        func_lut[191] = 204;  
        func_lut[192] = 204;  
        func_lut[193] = 203;  
        func_lut[194] = 203;  
        func_lut[195] = 203;  
        func_lut[196] = 202;  
        func_lut[197] = 202;  
        func_lut[198] = 202;  
        func_lut[199] = 202;  
        func_lut[200] = 201;  
        func_lut[201] = 201;  
        func_lut[202] = 201;  
        func_lut[203] = 200;  
        func_lut[204] = 200;  
        func_lut[205] = 200;  
        func_lut[206] = 200;  
        func_lut[207] = 199;  
        func_lut[208] = 199;  
        func_lut[209] = 199;  
        func_lut[210] = 199;  
        func_lut[211] = 198;  
        func_lut[212] = 198;  
        func_lut[213] = 198;  
        func_lut[214] = 197;  
        func_lut[215] = 197;  
        func_lut[216] = 197;  
        func_lut[217] = 197;  
        func_lut[218] = 196;  
        func_lut[219] = 196;  
        func_lut[220] = 196;  
        func_lut[221] = 196;  
        func_lut[222] = 195;  
        func_lut[223] = 195;  
        func_lut[224] = 195;  
        func_lut[225] = 195;  
        func_lut[226] = 194;  
        func_lut[227] = 194;  
        func_lut[228] = 194;  
        func_lut[229] = 193;  
        func_lut[230] = 193;  
        func_lut[231] = 193;  
        func_lut[232] = 193;  
        func_lut[233] = 192;  
        func_lut[234] = 192;  
        func_lut[235] = 192;  
        func_lut[236] = 192;  
        func_lut[237] = 191;  
        func_lut[238] = 191;  
        func_lut[239] = 191;  
        func_lut[240] = 191;  
        func_lut[241] = 190;  
        func_lut[242] = 190;  
        func_lut[243] = 190;  
        func_lut[244] = 190;  
        func_lut[245] = 189;  
        func_lut[246] = 189;  
        func_lut[247] = 189;  
        func_lut[248] = 189;  
        func_lut[249] = 188;  
        func_lut[250] = 188;  
        func_lut[251] = 188;  
        func_lut[252] = 188;  
        func_lut[253] = 187;  
        func_lut[254] = 187;  
        func_lut[255] = 187;  
        func_lut[256] = 187;  
        func_lut[257] = 186;  
        func_lut[258] = 186;  
        func_lut[259] = 186;  
        func_lut[260] = 186;  
        func_lut[261] = 185;  
        func_lut[262] = 185;  
        func_lut[263] = 185;  
        func_lut[264] = 185;  
        func_lut[265] = 184;  
        func_lut[266] = 184;  
        func_lut[267] = 184;  
        func_lut[268] = 184;  
        func_lut[269] = 183;  
        func_lut[270] = 183;  
        func_lut[271] = 183;  
        func_lut[272] = 183;  
        func_lut[273] = 182;  
        func_lut[274] = 182;  
        func_lut[275] = 182;  
        func_lut[276] = 182;  
        func_lut[277] = 182;  
        func_lut[278] = 181;  
        func_lut[279] = 181;  
        func_lut[280] = 181;  
        func_lut[281] = 181;  
        func_lut[282] = 180;  
        func_lut[283] = 180;  
        func_lut[284] = 180;  
        func_lut[285] = 180;  
        func_lut[286] = 179;  
        func_lut[287] = 179;  
        func_lut[288] = 179;  
        func_lut[289] = 179;  
        func_lut[290] = 178;  
        func_lut[291] = 178;  
        func_lut[292] = 178;  
        func_lut[293] = 178;  
        func_lut[294] = 178;  
        func_lut[295] = 177;  
        func_lut[296] = 177;  
        func_lut[297] = 177;  
        func_lut[298] = 177;  
        func_lut[299] = 176;  
        func_lut[300] = 176;  
        func_lut[301] = 176;  
        func_lut[302] = 176;  
        func_lut[303] = 175;  
        func_lut[304] = 175;  
        func_lut[305] = 175;  
        func_lut[306] = 175;  
        func_lut[307] = 175;  
        func_lut[308] = 174;  
        func_lut[309] = 174;  
        func_lut[310] = 174;  
        func_lut[311] = 174;  
        func_lut[312] = 173;  
        func_lut[313] = 173;  
        func_lut[314] = 173;  
        func_lut[315] = 173;  
        func_lut[316] = 173;  
        func_lut[317] = 172;  
        func_lut[318] = 172;  
        func_lut[319] = 172;  
        func_lut[320] = 172;  
        func_lut[321] = 171;  
        func_lut[322] = 171;  
        func_lut[323] = 171;  
        func_lut[324] = 171;  
        func_lut[325] = 171;  
        func_lut[326] = 170;  
        func_lut[327] = 170;  
        func_lut[328] = 170;  
        func_lut[329] = 170;  
        func_lut[330] = 170;  
        func_lut[331] = 169;  
        func_lut[332] = 169;  
        func_lut[333] = 169;  
        func_lut[334] = 169;  
        func_lut[335] = 168;  
        func_lut[336] = 168;  
        func_lut[337] = 168;  
        func_lut[338] = 168;  
        func_lut[339] = 168;  
        func_lut[340] = 167;  
        func_lut[341] = 167;  
        func_lut[342] = 167;  
        func_lut[343] = 167;  
        func_lut[344] = 167;  
        func_lut[345] = 166;  
        func_lut[346] = 166;  
        func_lut[347] = 166;  
        func_lut[348] = 166;  
        func_lut[349] = 166;  
        func_lut[350] = 165;  
        func_lut[351] = 165;  
        func_lut[352] = 165;  
        func_lut[353] = 165;  
        func_lut[354] = 165;  
        func_lut[355] = 164;  
        func_lut[356] = 164;  
        func_lut[357] = 164;  
        func_lut[358] = 164;  
        func_lut[359] = 163;  
        func_lut[360] = 163;  
        func_lut[361] = 163;  
        func_lut[362] = 163;  
        func_lut[363] = 163;  
        func_lut[364] = 162;  
        func_lut[365] = 162;  
        func_lut[366] = 162;  
        func_lut[367] = 162;  
        func_lut[368] = 162;  
        func_lut[369] = 161;  
        func_lut[370] = 161;  
        func_lut[371] = 161;  
        func_lut[372] = 161;  
        func_lut[373] = 161;  
        func_lut[374] = 160;  
        func_lut[375] = 160;  
        func_lut[376] = 160;  
        func_lut[377] = 160;  
        func_lut[378] = 160;  
        func_lut[379] = 160;  
        func_lut[380] = 159;  
        func_lut[381] = 159;  
        func_lut[382] = 159;  
        func_lut[383] = 159;  
        func_lut[384] = 159;  
        func_lut[385] = 158;  
        func_lut[386] = 158;  
        func_lut[387] = 158;  
        func_lut[388] = 158;  
        func_lut[389] = 158;  
        func_lut[390] = 157;  
        func_lut[391] = 157;  
        func_lut[392] = 157;  
        func_lut[393] = 157;  
        func_lut[394] = 157;  
        func_lut[395] = 156;  
        func_lut[396] = 156;  
        func_lut[397] = 156;  
        func_lut[398] = 156;  
        func_lut[399] = 156;  
        func_lut[400] = 155;  
        func_lut[401] = 155;  
        func_lut[402] = 155;  
        func_lut[403] = 155;  
        func_lut[404] = 155;  
        func_lut[405] = 155;  
        func_lut[406] = 154;  
        func_lut[407] = 154;  
        func_lut[408] = 154;  
        func_lut[409] = 154;  
        func_lut[410] = 154;  
        func_lut[411] = 153;  
        func_lut[412] = 153;  
        func_lut[413] = 153;  
        func_lut[414] = 153;  
        func_lut[415] = 153;  
        func_lut[416] = 153;  
        func_lut[417] = 152;  
        func_lut[418] = 152;  
        func_lut[419] = 152;  
        func_lut[420] = 152;  
        func_lut[421] = 152;  
        func_lut[422] = 151;  
        func_lut[423] = 151;  
        func_lut[424] = 151;  
        func_lut[425] = 151;  
        func_lut[426] = 151;  
        func_lut[427] = 151;  
        func_lut[428] = 150;  
        func_lut[429] = 150;  
        func_lut[430] = 150;  
        func_lut[431] = 150;  
        func_lut[432] = 150;  
        func_lut[433] = 149;  
        func_lut[434] = 149;  
        func_lut[435] = 149;  
        func_lut[436] = 149;  
        func_lut[437] = 149;  
        func_lut[438] = 149;  
        func_lut[439] = 148;  
        func_lut[440] = 148;  
        func_lut[441] = 148;  
        func_lut[442] = 148;  
        func_lut[443] = 148;  
        func_lut[444] = 148;  
        func_lut[445] = 147;  
        func_lut[446] = 147;  
        func_lut[447] = 147;  
        func_lut[448] = 147;  
        func_lut[449] = 147;  
        func_lut[450] = 146;  
        func_lut[451] = 146;  
        func_lut[452] = 146;  
        func_lut[453] = 146;  
        func_lut[454] = 146;  
        func_lut[455] = 146;  
        func_lut[456] = 145;  
        func_lut[457] = 145;  
        func_lut[458] = 145;  
        func_lut[459] = 145;  
        func_lut[460] = 145;  
        func_lut[461] = 145;  
        func_lut[462] = 144;  
        func_lut[463] = 144;  
        func_lut[464] = 144;  
        func_lut[465] = 144;  
        func_lut[466] = 144;  
        func_lut[467] = 144;  
        func_lut[468] = 143;  
        func_lut[469] = 143;  
        func_lut[470] = 143;  
        func_lut[471] = 143;  
        func_lut[472] = 143;  
        func_lut[473] = 143;  
        func_lut[474] = 142;  
        func_lut[475] = 142;  
        func_lut[476] = 142;  
        func_lut[477] = 142;  
        func_lut[478] = 142;  
        func_lut[479] = 142;  
        func_lut[480] = 141;  
        func_lut[481] = 141;  
        func_lut[482] = 141;  
        func_lut[483] = 141;  
        func_lut[484] = 141;  
        func_lut[485] = 141;  
        func_lut[486] = 140;  
        func_lut[487] = 140;  
        func_lut[488] = 140;  
        func_lut[489] = 140;  
        func_lut[490] = 140;  
        func_lut[491] = 140;  
        func_lut[492] = 140;  
        func_lut[493] = 139;  
        func_lut[494] = 139;  
        func_lut[495] = 139;  
        func_lut[496] = 139;  
        func_lut[497] = 139;  
        func_lut[498] = 139;  
        func_lut[499] = 138;  
        func_lut[500] = 138;  
        func_lut[501] = 138;  
        func_lut[502] = 138;  
        func_lut[503] = 138;  
        func_lut[504] = 138;  
        func_lut[505] = 137;  
        func_lut[506] = 137;  
        func_lut[507] = 137;  
        func_lut[508] = 137;  
        func_lut[509] = 137;  
        func_lut[510] = 137;  
        func_lut[511] = 137;  
        func_lut[512] = 136;  
        func_lut[513] = 136;  
        func_lut[514] = 136;  
        func_lut[515] = 136;  
        func_lut[516] = 136;  
        func_lut[517] = 136;  
        func_lut[518] = 135;  
        func_lut[519] = 135;  
        func_lut[520] = 135;  
        func_lut[521] = 135;  
        func_lut[522] = 135;  
        func_lut[523] = 135;  
        func_lut[524] = 135;  
        func_lut[525] = 134;  
        func_lut[526] = 134;  
        func_lut[527] = 134;  
        func_lut[528] = 134;  
        func_lut[529] = 134;  
        func_lut[530] = 134;  
        func_lut[531] = 133;  
        func_lut[532] = 133;  
        func_lut[533] = 133;  
        func_lut[534] = 133;  
        func_lut[535] = 133;  
        func_lut[536] = 133;  
        func_lut[537] = 133;  
        func_lut[538] = 132;  
        func_lut[539] = 132;  
        func_lut[540] = 132;  
        func_lut[541] = 132;  
        func_lut[542] = 132;  
        func_lut[543] = 132;  
        func_lut[544] = 132;  
        func_lut[545] = 131;  
        func_lut[546] = 131;  
        func_lut[547] = 131;  
        func_lut[548] = 131;  
        func_lut[549] = 131;  
        func_lut[550] = 131;  
        func_lut[551] = 131;  
        func_lut[552] = 130;  
        func_lut[553] = 130;  
        func_lut[554] = 130;  
        func_lut[555] = 130;  
        func_lut[556] = 130;  
        func_lut[557] = 130;  
        func_lut[558] = 130;  
        func_lut[559] = 129;  
        func_lut[560] = 129;  
        func_lut[561] = 129;  
        func_lut[562] = 129;  
        func_lut[563] = 129;  
        func_lut[564] = 129;  
        func_lut[565] = 129;  
        func_lut[566] = 128;  
        func_lut[567] = 128;  
        func_lut[568] = 128;  
        func_lut[569] = 128;  
        func_lut[570] = 128;  
        func_lut[571] = 128;  
        func_lut[572] = 128;  
        func_lut[573] = 127;  
        func_lut[574] = 127;  
        func_lut[575] = 127;  
        func_lut[576] = 127;  
        func_lut[577] = 127;  
        func_lut[578] = 127;  
        func_lut[579] = 127;  
        func_lut[580] = 126;  
        func_lut[581] = 126;  
        func_lut[582] = 126;  
        func_lut[583] = 126;  
        func_lut[584] = 126;  
        func_lut[585] = 126;  
        func_lut[586] = 126;  
        func_lut[587] = 125;  
        func_lut[588] = 125;  
        func_lut[589] = 125;  
        func_lut[590] = 125;  
        func_lut[591] = 125;  
        func_lut[592] = 125;  
        func_lut[593] = 125;  
        func_lut[594] = 125;  
        func_lut[595] = 124;  
        func_lut[596] = 124;  
        func_lut[597] = 124;  
        func_lut[598] = 124;  
        func_lut[599] = 124;  
        func_lut[600] = 124;  
        func_lut[601] = 124;  
        func_lut[602] = 123;  
        func_lut[603] = 123;  
        func_lut[604] = 123;  
        func_lut[605] = 123;  
        func_lut[606] = 123;  
        func_lut[607] = 123;  
        func_lut[608] = 123;  
        func_lut[609] = 123;  
        func_lut[610] = 122;  
        func_lut[611] = 122;  
        func_lut[612] = 122;  
        func_lut[613] = 122;  
        func_lut[614] = 122;  
        func_lut[615] = 122;  
        func_lut[616] = 122;  
        func_lut[617] = 121;  
        func_lut[618] = 121;  
        func_lut[619] = 121;  
        func_lut[620] = 121;  
        func_lut[621] = 121;  
        func_lut[622] = 121;  
        func_lut[623] = 121;  
        func_lut[624] = 121;  
        func_lut[625] = 120;  
        func_lut[626] = 120;  
        func_lut[627] = 120;  
        func_lut[628] = 120;  
        func_lut[629] = 120;  
        func_lut[630] = 120;  
        func_lut[631] = 120;  
        func_lut[632] = 120;  
        func_lut[633] = 119;  
        func_lut[634] = 119;  
        func_lut[635] = 119;  
        func_lut[636] = 119;  
        func_lut[637] = 119;  
        func_lut[638] = 119;  
        func_lut[639] = 119;  
        func_lut[640] = 119;  
        func_lut[641] = 118;  
        func_lut[642] = 118;  
        func_lut[643] = 118;  
        func_lut[644] = 118;  
        func_lut[645] = 118;  
        func_lut[646] = 118;  
        func_lut[647] = 118;  
        func_lut[648] = 118;  
        func_lut[649] = 117;  
        func_lut[650] = 117;  
        func_lut[651] = 117;  
        func_lut[652] = 117;  
        func_lut[653] = 117;  
        func_lut[654] = 117;  
        func_lut[655] = 117;  
        func_lut[656] = 117;  
        func_lut[657] = 116;  
        func_lut[658] = 116;  
        func_lut[659] = 116;  
        func_lut[660] = 116;  
        func_lut[661] = 116;  
        func_lut[662] = 116;  
        func_lut[663] = 116;  
        func_lut[664] = 116;  
        func_lut[665] = 115;  
        func_lut[666] = 115;  
        func_lut[667] = 115;  
        func_lut[668] = 115;  
        func_lut[669] = 115;  
        func_lut[670] = 115;  
        func_lut[671] = 115;  
        func_lut[672] = 115;  
        func_lut[673] = 115;  
        func_lut[674] = 114;  
        func_lut[675] = 114;  
        func_lut[676] = 114;  
        func_lut[677] = 114;  
        func_lut[678] = 114;  
        func_lut[679] = 114;  
        func_lut[680] = 114;  
        func_lut[681] = 114;  
        func_lut[682] = 113;  
        func_lut[683] = 113;  
        func_lut[684] = 113;  
        func_lut[685] = 113;  
        func_lut[686] = 113;  
        func_lut[687] = 113;  
        func_lut[688] = 113;  
        func_lut[689] = 113;  
        func_lut[690] = 113;  
        func_lut[691] = 112;  
        func_lut[692] = 112;  
        func_lut[693] = 112;  
        func_lut[694] = 112;  
        func_lut[695] = 112;  
        func_lut[696] = 112;  
        func_lut[697] = 112;  
        func_lut[698] = 112;  
        func_lut[699] = 111;  
        func_lut[700] = 111;  
        func_lut[701] = 111;  
        func_lut[702] = 111;  
        func_lut[703] = 111;  
        func_lut[704] = 111;  
        func_lut[705] = 111;  
        func_lut[706] = 111;  
        func_lut[707] = 111;  
        func_lut[708] = 110;  
        func_lut[709] = 110;  
        func_lut[710] = 110;  
        func_lut[711] = 110;  
        func_lut[712] = 110;  
        func_lut[713] = 110;  
        func_lut[714] = 110;  
        func_lut[715] = 110;  
        func_lut[716] = 110;  
        func_lut[717] = 109;  
        func_lut[718] = 109;  
        func_lut[719] = 109;  
        func_lut[720] = 109;  
        func_lut[721] = 109;  
        func_lut[722] = 109;  
        func_lut[723] = 109;  
        func_lut[724] = 109;  
        func_lut[725] = 109;  
        func_lut[726] = 108;  
        func_lut[727] = 108;  
        func_lut[728] = 108;  
        func_lut[729] = 108;  
        func_lut[730] = 108;  
        func_lut[731] = 108;  
        func_lut[732] = 108;  
        func_lut[733] = 108;  
        func_lut[734] = 108;  
        func_lut[735] = 107;  
        func_lut[736] = 107;  
        func_lut[737] = 107;  
        func_lut[738] = 107;  
        func_lut[739] = 107;  
        func_lut[740] = 107;  
        func_lut[741] = 107;  
        func_lut[742] = 107;  
        func_lut[743] = 107;  
        func_lut[744] = 107;  
        func_lut[745] = 106;  
        func_lut[746] = 106;  
        func_lut[747] = 106;  
        func_lut[748] = 106;  
        func_lut[749] = 106;  
        func_lut[750] = 106;  
        func_lut[751] = 106;  
        func_lut[752] = 106;  
        func_lut[753] = 106;  
        func_lut[754] = 105;  
        func_lut[755] = 105;  
        func_lut[756] = 105;  
        func_lut[757] = 105;  
        func_lut[758] = 105;  
        func_lut[759] = 105;  
        func_lut[760] = 105;  
        func_lut[761] = 105;  
        func_lut[762] = 105;  
        func_lut[763] = 105;  
        func_lut[764] = 104;  
        func_lut[765] = 104;  
        func_lut[766] = 104;  
        func_lut[767] = 104;  
        func_lut[768] = 104;  
        func_lut[769] = 104;  
        func_lut[770] = 104;  
        func_lut[771] = 104;  
        func_lut[772] = 104;  
        func_lut[773] = 103;  
        func_lut[774] = 103;  
        func_lut[775] = 103;  
        func_lut[776] = 103;  
        func_lut[777] = 103;  
        func_lut[778] = 103;  
        func_lut[779] = 103;  
        func_lut[780] = 103;  
        func_lut[781] = 103;  
        func_lut[782] = 103;  
        func_lut[783] = 102;  
        func_lut[784] = 102;  
        func_lut[785] = 102;  
        func_lut[786] = 102;  
        func_lut[787] = 102;  
        func_lut[788] = 102;  
        func_lut[789] = 102;  
        func_lut[790] = 102;  
        func_lut[791] = 102;  
        func_lut[792] = 102;  
        func_lut[793] = 101;  
        func_lut[794] = 101;  
        func_lut[795] = 101;  
        func_lut[796] = 101;  
        func_lut[797] = 101;  
        func_lut[798] = 101;  
        func_lut[799] = 101;  
        func_lut[800] = 101;  
        func_lut[801] = 101;  
        func_lut[802] = 101;  
        func_lut[803] = 100;  
        func_lut[804] = 100;  
        func_lut[805] = 100;  
        func_lut[806] = 100;  
        func_lut[807] = 100;  
        func_lut[808] = 100;  
        func_lut[809] = 100;  
        func_lut[810] = 100;  
        func_lut[811] = 100;  
        func_lut[812] = 100;  
        func_lut[813] = 100;  
        func_lut[814] = 99;  
        func_lut[815] = 99;  
        func_lut[816] = 99;  
        func_lut[817] = 99;  
        func_lut[818] = 99;  
        func_lut[819] = 99;  
        func_lut[820] = 99;  
        func_lut[821] = 99;  
        func_lut[822] = 99;  
        func_lut[823] = 99;  
        func_lut[824] = 98;  
        func_lut[825] = 98;  
        func_lut[826] = 98;  
        func_lut[827] = 98;  
        func_lut[828] = 98;  
        func_lut[829] = 98;  
        func_lut[830] = 98;  
        func_lut[831] = 98;  
        func_lut[832] = 98;  
        func_lut[833] = 98;  
        func_lut[834] = 98;  
        func_lut[835] = 97;  
        func_lut[836] = 97;  
        func_lut[837] = 97;  
        func_lut[838] = 97;  
        func_lut[839] = 97;  
        func_lut[840] = 97;  
        func_lut[841] = 97;  
        func_lut[842] = 97;  
        func_lut[843] = 97;  
        func_lut[844] = 97;  
        func_lut[845] = 96;  
        func_lut[846] = 96;  
        func_lut[847] = 96;  
        func_lut[848] = 96;  
        func_lut[849] = 96;  
        func_lut[850] = 96;  
        func_lut[851] = 96;  
        func_lut[852] = 96;  
        func_lut[853] = 96;  
        func_lut[854] = 96;  
        func_lut[855] = 96;  
        func_lut[856] = 95;  
        func_lut[857] = 95;  
        func_lut[858] = 95;  
        func_lut[859] = 95;  
        func_lut[860] = 95;  
        func_lut[861] = 95;  
        func_lut[862] = 95;  
        func_lut[863] = 95;  
        func_lut[864] = 95;  
        func_lut[865] = 95;  
        func_lut[866] = 95;  
        func_lut[867] = 94;  
        func_lut[868] = 94;  
        func_lut[869] = 94;  
        func_lut[870] = 94;  
        func_lut[871] = 94;  
        func_lut[872] = 94;  
        func_lut[873] = 94;  
        func_lut[874] = 94;  
        func_lut[875] = 94;  
        func_lut[876] = 94;  
        func_lut[877] = 94;  
        func_lut[878] = 94;  
        func_lut[879] = 93;  
        func_lut[880] = 93;  
        func_lut[881] = 93;  
        func_lut[882] = 93;  
        func_lut[883] = 93;  
        func_lut[884] = 93;  
        func_lut[885] = 93;  
        func_lut[886] = 93;  
        func_lut[887] = 93;  
        func_lut[888] = 93;  
        func_lut[889] = 93;  
        func_lut[890] = 92;  
        func_lut[891] = 92;  
        func_lut[892] = 92;  
        func_lut[893] = 92;  
        func_lut[894] = 92;  
        func_lut[895] = 92;  
        func_lut[896] = 92;  
        func_lut[897] = 92;  
        func_lut[898] = 92;  
        func_lut[899] = 92;  
        func_lut[900] = 92;  
        func_lut[901] = 92;  
        func_lut[902] = 91;  
        func_lut[903] = 91;  
        func_lut[904] = 91;  
        func_lut[905] = 91;  
        func_lut[906] = 91;  
        func_lut[907] = 91;  
        func_lut[908] = 91;  
        func_lut[909] = 91;  
        func_lut[910] = 91;  
        func_lut[911] = 91;  
        func_lut[912] = 91;  
        func_lut[913] = 91;  
        func_lut[914] = 90;  
        func_lut[915] = 90;  
        func_lut[916] = 90;  
        func_lut[917] = 90;  
        func_lut[918] = 90;  
        func_lut[919] = 90;  
        func_lut[920] = 90;  
        func_lut[921] = 90;  
        func_lut[922] = 90;  
        func_lut[923] = 90;  
        func_lut[924] = 90;  
        func_lut[925] = 90;  
        func_lut[926] = 89;  
        func_lut[927] = 89;  
        func_lut[928] = 89;  
        func_lut[929] = 89;  
        func_lut[930] = 89;  
        func_lut[931] = 89;  
        func_lut[932] = 89;  
        func_lut[933] = 89;  
        func_lut[934] = 89;  
        func_lut[935] = 89;  
        func_lut[936] = 89;  
        func_lut[937] = 89;  
        func_lut[938] = 88;  
        func_lut[939] = 88;  
        func_lut[940] = 88;  
        func_lut[941] = 88;  
        func_lut[942] = 88;  
        func_lut[943] = 88;  
        func_lut[944] = 88;  
        func_lut[945] = 88;  
        func_lut[946] = 88;  
        func_lut[947] = 88;  
        func_lut[948] = 88;  
        func_lut[949] = 88;  
        func_lut[950] = 88;  
        func_lut[951] = 87;  
        func_lut[952] = 87;  
        func_lut[953] = 87;  
        func_lut[954] = 87;  
        func_lut[955] = 87;  
        func_lut[956] = 87;  
        func_lut[957] = 87;  
        func_lut[958] = 87;  
        func_lut[959] = 87;  
        func_lut[960] = 87;  
        func_lut[961] = 87;  
        func_lut[962] = 87;  
        func_lut[963] = 86;  
        func_lut[964] = 86;  
        func_lut[965] = 86;  
        func_lut[966] = 86;  
        func_lut[967] = 86;  
        func_lut[968] = 86;  
        func_lut[969] = 86;  
        func_lut[970] = 86;  
        func_lut[971] = 86;  
        func_lut[972] = 86;  
        func_lut[973] = 86;  
        func_lut[974] = 86;  
        func_lut[975] = 86;  
        func_lut[976] = 85;  
        func_lut[977] = 85;  
        func_lut[978] = 85;  
        func_lut[979] = 85;  
        func_lut[980] = 85;  
        func_lut[981] = 85;  
        func_lut[982] = 85;  
        func_lut[983] = 85;  
        func_lut[984] = 85;  
        func_lut[985] = 85;  
        func_lut[986] = 85;  
        func_lut[987] = 85;  
        func_lut[988] = 85;  
        func_lut[989] = 84;  
        func_lut[990] = 84;  
        func_lut[991] = 84;  
        func_lut[992] = 84;  
        func_lut[993] = 84;  
        func_lut[994] = 84;  
        func_lut[995] = 84;  
        func_lut[996] = 84;  
        func_lut[997] = 84;  
        func_lut[998] = 84;  
        func_lut[999] = 84;  
        func_lut[1000] = 84;  
        func_lut[1001] = 84;  
        func_lut[1002] = 84;  
        func_lut[1003] = 83;  
        func_lut[1004] = 83;  
        func_lut[1005] = 83;  
        func_lut[1006] = 83;  
        func_lut[1007] = 83;  
        func_lut[1008] = 83;  
        func_lut[1009] = 83;  
        func_lut[1010] = 83;  
        func_lut[1011] = 83;  
        func_lut[1012] = 83;  
        func_lut[1013] = 83;  
        func_lut[1014] = 83;  
        func_lut[1015] = 83;  
        func_lut[1016] = 82;  
        func_lut[1017] = 82;  
        func_lut[1018] = 82;  
        func_lut[1019] = 82;  
        func_lut[1020] = 82;  
        func_lut[1021] = 82;  
        func_lut[1022] = 82;  
        func_lut[1023] = 82;  
        func_lut[1024] = 8179;  
        func_lut[1025] = 8107;  
        func_lut[1026] = 8037;  
        func_lut[1027] = 7968;  
        func_lut[1028] = 7899;  
        func_lut[1029] = 7831;  
        func_lut[1030] = 7764;  
        func_lut[1031] = 7698;  
        func_lut[1032] = 7633;  
        func_lut[1033] = 7569;  
        func_lut[1034] = 7505;  
        func_lut[1035] = 7443;  
        func_lut[1036] = 7381;  
        func_lut[1037] = 7319;  
        func_lut[1038] = 7259;  
        func_lut[1039] = 7199;  
        func_lut[1040] = 7140;  
        func_lut[1041] = 7082;  
        func_lut[1042] = 7025;  
        func_lut[1043] = 6968;  
        func_lut[1044] = 6912;  
        func_lut[1045] = 6856;  
        func_lut[1046] = 6801;  
        func_lut[1047] = 6747;  
        func_lut[1048] = 6694;  
        func_lut[1049] = 6641;  
        func_lut[1050] = 6589;  
        func_lut[1051] = 6537;  
        func_lut[1052] = 6486;  
        func_lut[1053] = 6436;  
        func_lut[1054] = 6386;  
        func_lut[1055] = 6336;  
        func_lut[1056] = 6288;  
        func_lut[1057] = 6240;  
        func_lut[1058] = 6192;  
        func_lut[1059] = 6145;  
        func_lut[1060] = 6098;  
        func_lut[1061] = 6052;  
        func_lut[1062] = 6007;  
        func_lut[1063] = 5962;  
        func_lut[1064] = 5918;  
        func_lut[1065] = 5874;  
        func_lut[1066] = 5830;  
        func_lut[1067] = 5787;  
        func_lut[1068] = 5745;  
        func_lut[1069] = 5703;  
        func_lut[1070] = 5661;  
        func_lut[1071] = 5620;  
        func_lut[1072] = 5579;  
        func_lut[1073] = 5539;  
        func_lut[1074] = 5499;  
        func_lut[1075] = 5460;  
        func_lut[1076] = 5421;  
        func_lut[1077] = 5382;  
        func_lut[1078] = 5344;  
        func_lut[1079] = 5306;  
        func_lut[1080] = 5269;  
        func_lut[1081] = 5232;  
        func_lut[1082] = 5195;  
        func_lut[1083] = 5159;  
        func_lut[1084] = 5124;  
        func_lut[1085] = 5088;  
        func_lut[1086] = 5053;  
        func_lut[1087] = 5018;  
        func_lut[1088] = 4984;  
        func_lut[1089] = 4950;  
        func_lut[1090] = 4916;  
        func_lut[1091] = 4883;  
        func_lut[1092] = 4850;  
        func_lut[1093] = 4817;  
        func_lut[1094] = 4785;  
        func_lut[1095] = 4753;  
        func_lut[1096] = 4721;  
        func_lut[1097] = 4690;  
        func_lut[1098] = 4659;  
        func_lut[1099] = 4628;  
        func_lut[1100] = 4598;  
        func_lut[1101] = 4568;  
        func_lut[1102] = 4538;  
        func_lut[1103] = 4508;  
        func_lut[1104] = 4479;  
        func_lut[1105] = 4450;  
        func_lut[1106] = 4422;  
        func_lut[1107] = 4393;  
        func_lut[1108] = 4365;  
        func_lut[1109] = 4337;  
        func_lut[1110] = 4310;  
        func_lut[1111] = 4282;  
        func_lut[1112] = 4255;  
        func_lut[1113] = 4228;  
        func_lut[1114] = 4202;  
        func_lut[1115] = 4175;  
        func_lut[1116] = 4149;  
        func_lut[1117] = 4123;  
        func_lut[1118] = 4098;  
        func_lut[1119] = 4073;  
        func_lut[1120] = 4047;  
        func_lut[1121] = 4023;  
        func_lut[1122] = 3998;  
        func_lut[1123] = 3973;  
        func_lut[1124] = 3949;  
        func_lut[1125] = 3925;  
        func_lut[1126] = 3901;  
        func_lut[1127] = 3878;  
        func_lut[1128] = 3855;  
        func_lut[1129] = 3831;  
        func_lut[1130] = 3808;  
        func_lut[1131] = 3786;  
        func_lut[1132] = 3763;  
        func_lut[1133] = 3741;  
        func_lut[1134] = 3719;  
        func_lut[1135] = 3697;  
        func_lut[1136] = 3675;  
        func_lut[1137] = 3654;  
        func_lut[1138] = 3632;  
        func_lut[1139] = 3611;  
        func_lut[1140] = 3590;  
        func_lut[1141] = 3569;  
        func_lut[1142] = 3549;  
        func_lut[1143] = 3528;  
        func_lut[1144] = 3508;  
        func_lut[1145] = 3488;  
        func_lut[1146] = 3468;  
        func_lut[1147] = 3448;  
        func_lut[1148] = 3429;  
        func_lut[1149] = 3409;  
        func_lut[1150] = 3390;  
        func_lut[1151] = 3371;  
        func_lut[1152] = 3352;  
        func_lut[1153] = 3333;  
        func_lut[1154] = 3315;  
        func_lut[1155] = 3296;  
        func_lut[1156] = 3278;  
        func_lut[1157] = 3260;  
        func_lut[1158] = 3242;  
        func_lut[1159] = 3224;  
        func_lut[1160] = 3206;  
        func_lut[1161] = 3189;  
        func_lut[1162] = 3171;  
        func_lut[1163] = 3154;  
        func_lut[1164] = 3137;  
        func_lut[1165] = 3120;  
        func_lut[1166] = 3103;  
        func_lut[1167] = 3086;  
        func_lut[1168] = 3070;  
        func_lut[1169] = 3053;  
        func_lut[1170] = 3037;  
        func_lut[1171] = 3021;  
        func_lut[1172] = 3005;  
        func_lut[1173] = 2989;  
        func_lut[1174] = 2973;  
        func_lut[1175] = 2957;  
        func_lut[1176] = 2942;  
        func_lut[1177] = 2926;  
        func_lut[1178] = 2911;  
        func_lut[1179] = 2896;  
        func_lut[1180] = 2881;  
        func_lut[1181] = 2866;  
        func_lut[1182] = 2851;  
        func_lut[1183] = 2836;  
        func_lut[1184] = 2822;  
        func_lut[1185] = 2807;  
        func_lut[1186] = 2793;  
        func_lut[1187] = 2778;  
        func_lut[1188] = 2764;  
        func_lut[1189] = 2750;  
        func_lut[1190] = 2736;  
        func_lut[1191] = 2722;  
        func_lut[1192] = 2709;  
        func_lut[1193] = 2695;  
        func_lut[1194] = 2681;  
        func_lut[1195] = 2668;  
        func_lut[1196] = 2655;  
        func_lut[1197] = 2641;  
        func_lut[1198] = 2628;  
        func_lut[1199] = 2615;  
        func_lut[1200] = 2602;  
        func_lut[1201] = 2589;  
        func_lut[1202] = 2577;  
        func_lut[1203] = 2564;  
        func_lut[1204] = 2552;  
        func_lut[1205] = 2539;  
        func_lut[1206] = 2527;  
        func_lut[1207] = 2514;  
        func_lut[1208] = 2502;  
        func_lut[1209] = 2490;  
        func_lut[1210] = 2478;  
        func_lut[1211] = 2466;  
        func_lut[1212] = 2454;  
        func_lut[1213] = 2443;  
        func_lut[1214] = 2431;  
        func_lut[1215] = 2419;  
        func_lut[1216] = 2408;  
        func_lut[1217] = 2396;  
        func_lut[1218] = 2385;  
        func_lut[1219] = 2374;  
        func_lut[1220] = 2362;  
        func_lut[1221] = 2351;  
        func_lut[1222] = 2340;  
        func_lut[1223] = 2329;  
        func_lut[1224] = 2319;  
        func_lut[1225] = 2308;  
        func_lut[1226] = 2297;  
        func_lut[1227] = 2286;  
        func_lut[1228] = 2276;  
        func_lut[1229] = 2265;  
        func_lut[1230] = 2255;  
        func_lut[1231] = 2244;  
        func_lut[1232] = 2234;  
        func_lut[1233] = 2224;  
        func_lut[1234] = 2214;  
        func_lut[1235] = 2204;  
        func_lut[1236] = 2194;  
        func_lut[1237] = 2184;  
        func_lut[1238] = 2174;  
        func_lut[1239] = 2164;  
        func_lut[1240] = 2154;  
        func_lut[1241] = 2145;  
        func_lut[1242] = 2135;  
        func_lut[1243] = 2125;  
        func_lut[1244] = 2116;  
        func_lut[1245] = 2107;  
        func_lut[1246] = 2097;  
        func_lut[1247] = 2088;  
        func_lut[1248] = 2079;  
        func_lut[1249] = 2070;  
        func_lut[1250] = 2060;  
        func_lut[1251] = 2051;  
        func_lut[1252] = 2042;  
        func_lut[1253] = 2033;  
        func_lut[1254] = 2025;  
        func_lut[1255] = 2016;  
        func_lut[1256] = 2007;  
        func_lut[1257] = 1998;  
        func_lut[1258] = 1990;  
        func_lut[1259] = 1981;  
        func_lut[1260] = 1973;  
        func_lut[1261] = 1964;  
        func_lut[1262] = 1956;  
        func_lut[1263] = 1947;  
        func_lut[1264] = 1939;  
        func_lut[1265] = 1931;  
        func_lut[1266] = 1922;  
        func_lut[1267] = 1914;  
        func_lut[1268] = 1906;  
        func_lut[1269] = 1898;  
        func_lut[1270] = 1890;  
        func_lut[1271] = 1882;  
        func_lut[1272] = 1874;  
        func_lut[1273] = 1866;  
        func_lut[1274] = 1859;  
        func_lut[1275] = 1851;  
        func_lut[1276] = 1843;  
        func_lut[1277] = 1835;  
        func_lut[1278] = 1828;  
        func_lut[1279] = 1820;  
        func_lut[1280] = 1813;  
        func_lut[1281] = 1805;  
        func_lut[1282] = 1798;  
        func_lut[1283] = 1790;  
        func_lut[1284] = 1783;  
        func_lut[1285] = 1776;  
        func_lut[1286] = 1769;  
        func_lut[1287] = 1761;  
        func_lut[1288] = 1754;  
        func_lut[1289] = 1747;  
        func_lut[1290] = 1740;  
        func_lut[1291] = 1733;  
        func_lut[1292] = 1726;  
        func_lut[1293] = 1719;  
        func_lut[1294] = 1712;  
        func_lut[1295] = 1705;  
        func_lut[1296] = 1699;  
        func_lut[1297] = 1692;  
        func_lut[1298] = 1685;  
        func_lut[1299] = 1678;  
        func_lut[1300] = 1672;  
        func_lut[1301] = 1665;  
        func_lut[1302] = 1658;  
        func_lut[1303] = 1652;  
        func_lut[1304] = 1645;  
        func_lut[1305] = 1639;  
        func_lut[1306] = 1633;  
        func_lut[1307] = 1626;  
        func_lut[1308] = 1620;  
        func_lut[1309] = 1614;  
        func_lut[1310] = 1607;  
        func_lut[1311] = 1601;  
        func_lut[1312] = 1595;  
        func_lut[1313] = 1589;  
        func_lut[1314] = 1582;  
        func_lut[1315] = 1576;  
        func_lut[1316] = 1570;  
        func_lut[1317] = 1564;  
        func_lut[1318] = 1558;  
        func_lut[1319] = 1552;  
        func_lut[1320] = 1546;  
        func_lut[1321] = 1541;  
        func_lut[1322] = 1535;  
        func_lut[1323] = 1529;  
        func_lut[1324] = 1523;  
        func_lut[1325] = 1517;  
        func_lut[1326] = 1512;  
        func_lut[1327] = 1506;  
        func_lut[1328] = 1500;  
        func_lut[1329] = 1495;  
        func_lut[1330] = 1489;  
        func_lut[1331] = 1483;  
        func_lut[1332] = 1478;  
        func_lut[1333] = 1472;  
        func_lut[1334] = 1467;  
        func_lut[1335] = 1462;  
        func_lut[1336] = 1456;  
        func_lut[1337] = 1451;  
        func_lut[1338] = 1445;  
        func_lut[1339] = 1440;  
        func_lut[1340] = 1435;  
        func_lut[1341] = 1430;  
        func_lut[1342] = 1424;  
        func_lut[1343] = 1419;  
        func_lut[1344] = 1414;  
        func_lut[1345] = 1409;  
        func_lut[1346] = 1404;  
        func_lut[1347] = 1399;  
        func_lut[1348] = 1393;  
        func_lut[1349] = 1388;  
        func_lut[1350] = 1383;  
        func_lut[1351] = 1378;  
        func_lut[1352] = 1373;  
        func_lut[1353] = 1369;  
        func_lut[1354] = 1364;  
        func_lut[1355] = 1359;  
        func_lut[1356] = 1354;  
        func_lut[1357] = 1349;  
        func_lut[1358] = 1344;  
        func_lut[1359] = 1340;  
        func_lut[1360] = 1335;  
        func_lut[1361] = 1330;  
        func_lut[1362] = 1325;  
        func_lut[1363] = 1321;  
        func_lut[1364] = 1316;  
        func_lut[1365] = 1311;  
        func_lut[1366] = 1307;  
        func_lut[1367] = 1302;  
        func_lut[1368] = 1298;  
        func_lut[1369] = 1293;  
        func_lut[1370] = 1289;  
        func_lut[1371] = 1284;  
        func_lut[1372] = 1280;  
        func_lut[1373] = 1275;  
        func_lut[1374] = 1271;  
        func_lut[1375] = 1266;  
        func_lut[1376] = 1262;  
        func_lut[1377] = 1258;  
        func_lut[1378] = 1253;  
        func_lut[1379] = 1249;  
        func_lut[1380] = 1245;  
        func_lut[1381] = 1241;  
        func_lut[1382] = 1236;  
        func_lut[1383] = 1232;  
        func_lut[1384] = 1228;  
        func_lut[1385] = 1224;  
        func_lut[1386] = 1220;  
        func_lut[1387] = 1216;  
        func_lut[1388] = 1211;  
        func_lut[1389] = 1207;  
        func_lut[1390] = 1203;  
        func_lut[1391] = 1199;  
        func_lut[1392] = 1195;  
        func_lut[1393] = 1191;  
        func_lut[1394] = 1187;  
        func_lut[1395] = 1183;  
        func_lut[1396] = 1179;  
        func_lut[1397] = 1175;  
        func_lut[1398] = 1172;  
        func_lut[1399] = 1168;  
        func_lut[1400] = 1164;  
        func_lut[1401] = 1160;  
        func_lut[1402] = 1156;  
        func_lut[1403] = 1152;  
        func_lut[1404] = 1148;  
        func_lut[1405] = 1145;  
        func_lut[1406] = 1141;  
        func_lut[1407] = 1137;  
        func_lut[1408] = 1134;  
        func_lut[1409] = 1130;  
        func_lut[1410] = 1126;  
        func_lut[1411] = 1122;  
        func_lut[1412] = 1119;  
        func_lut[1413] = 1115;  
        func_lut[1414] = 1112;  
        func_lut[1415] = 1108;  
        func_lut[1416] = 1104;  
        func_lut[1417] = 1101;  
        func_lut[1418] = 1097;  
        func_lut[1419] = 1094;  
        func_lut[1420] = 1090;  
        func_lut[1421] = 1087;  
        func_lut[1422] = 1083;  
        func_lut[1423] = 1080;  
        func_lut[1424] = 1076;  
        func_lut[1425] = 1073;  
        func_lut[1426] = 1070;  
        func_lut[1427] = 1066;  
        func_lut[1428] = 1063;  
        func_lut[1429] = 1060;  
        func_lut[1430] = 1056;  
        func_lut[1431] = 1053;  
        func_lut[1432] = 1050;  
        func_lut[1433] = 1046;  
        func_lut[1434] = 1043;  
        func_lut[1435] = 1040;  
        func_lut[1436] = 1036;  
        func_lut[1437] = 1033;  
        func_lut[1438] = 1030;  
        func_lut[1439] = 1027;  
        func_lut[1440] = 1024;  
        func_lut[1441] = 1020;  
        func_lut[1442] = 1017;  
        func_lut[1443] = 1014;  
        func_lut[1444] = 1011;  
        func_lut[1445] = 1008;  
        func_lut[1446] = 1005;  
        func_lut[1447] = 1002;  
        func_lut[1448] = 999;  
        func_lut[1449] = 996;  
        func_lut[1450] = 993;  
        func_lut[1451] = 990;  
        func_lut[1452] = 987;  
        func_lut[1453] = 984;  
        func_lut[1454] = 981;  
        func_lut[1455] = 978;  
        func_lut[1456] = 975;  
        func_lut[1457] = 972;  
        func_lut[1458] = 969;  
        func_lut[1459] = 966;  
        func_lut[1460] = 963;  
        func_lut[1461] = 960;  
        func_lut[1462] = 957;  
        func_lut[1463] = 954;  
        func_lut[1464] = 951;  
        func_lut[1465] = 949;  
        func_lut[1466] = 946;  
        func_lut[1467] = 943;  
        func_lut[1468] = 940;  
        func_lut[1469] = 937;  
        func_lut[1470] = 935;  
        func_lut[1471] = 932;  
        func_lut[1472] = 929;  
        func_lut[1473] = 926;  
        func_lut[1474] = 924;  
        func_lut[1475] = 921;  
        func_lut[1476] = 918;  
        func_lut[1477] = 915;  
        func_lut[1478] = 913;  
        func_lut[1479] = 910;  
        func_lut[1480] = 907;  
        func_lut[1481] = 905;  
        func_lut[1482] = 902;  
        func_lut[1483] = 899;  
        func_lut[1484] = 897;  
        func_lut[1485] = 894;  
        func_lut[1486] = 892;  
        func_lut[1487] = 889;  
        func_lut[1488] = 887;  
        func_lut[1489] = 884;  
        func_lut[1490] = 881;  
        func_lut[1491] = 879;  
        func_lut[1492] = 876;  
        func_lut[1493] = 874;  
        func_lut[1494] = 871;  
        func_lut[1495] = 869;  
        func_lut[1496] = 866;  
        func_lut[1497] = 864;  
        func_lut[1498] = 861;  
        func_lut[1499] = 859;  
        func_lut[1500] = 857;  
        func_lut[1501] = 854;  
        func_lut[1502] = 852;  
        func_lut[1503] = 849;  
        func_lut[1504] = 847;  
        func_lut[1505] = 844;  
        func_lut[1506] = 842;  
        func_lut[1507] = 840;  
        func_lut[1508] = 837;  
        func_lut[1509] = 835;  
        func_lut[1510] = 833;  
        func_lut[1511] = 830;  
        func_lut[1512] = 828;  
        func_lut[1513] = 826;  
        func_lut[1514] = 823;  
        func_lut[1515] = 821;  
        func_lut[1516] = 819;  
        func_lut[1517] = 817;  
        func_lut[1518] = 814;  
        func_lut[1519] = 812;  
        func_lut[1520] = 810;  
        func_lut[1521] = 808;  
        func_lut[1522] = 805;  
        func_lut[1523] = 803;  
        func_lut[1524] = 801;  
        func_lut[1525] = 799;  
        func_lut[1526] = 797;  
        func_lut[1527] = 794;  
        func_lut[1528] = 792;  
        func_lut[1529] = 790;  
        func_lut[1530] = 788;  
        func_lut[1531] = 786;  
        func_lut[1532] = 784;  
        func_lut[1533] = 782;  
        func_lut[1534] = 779;  
        func_lut[1535] = 777;  
        func_lut[1536] = 775;  
        func_lut[1537] = 773;  
        func_lut[1538] = 771;  
        func_lut[1539] = 769;  
        func_lut[1540] = 767;  
        func_lut[1541] = 765;  
        func_lut[1542] = 763;  
        func_lut[1543] = 761;  
        func_lut[1544] = 759;  
        func_lut[1545] = 757;  
        func_lut[1546] = 755;  
        func_lut[1547] = 753;  
        func_lut[1548] = 751;  
        func_lut[1549] = 749;  
        func_lut[1550] = 747;  
        func_lut[1551] = 745;  
        func_lut[1552] = 743;  
        func_lut[1553] = 741;  
        func_lut[1554] = 739;  
        func_lut[1555] = 737;  
        func_lut[1556] = 735;  
        func_lut[1557] = 733;  
        func_lut[1558] = 731;  
        func_lut[1559] = 729;  
        func_lut[1560] = 727;  
        func_lut[1561] = 725;  
        func_lut[1562] = 723;  
        func_lut[1563] = 722;  
        func_lut[1564] = 720;  
        func_lut[1565] = 718;  
        func_lut[1566] = 716;  
        func_lut[1567] = 714;  
        func_lut[1568] = 712;  
        func_lut[1569] = 710;  
        func_lut[1570] = 709;  
        func_lut[1571] = 707;  
        func_lut[1572] = 705;  
        func_lut[1573] = 703;  
        func_lut[1574] = 701;  
        func_lut[1575] = 699;  
        func_lut[1576] = 698;  
        func_lut[1577] = 696;  
        func_lut[1578] = 694;  
        func_lut[1579] = 692;  
        func_lut[1580] = 691;  
        func_lut[1581] = 689;  
        func_lut[1582] = 687;  
        func_lut[1583] = 685;  
        func_lut[1584] = 684;  
        func_lut[1585] = 682;  
        func_lut[1586] = 680;  
        func_lut[1587] = 678;  
        func_lut[1588] = 677;  
        func_lut[1589] = 675;  
        func_lut[1590] = 673;  
        func_lut[1591] = 672;  
        func_lut[1592] = 670;  
        func_lut[1593] = 668;  
        func_lut[1594] = 667;  
        func_lut[1595] = 665;  
        func_lut[1596] = 663;  
        func_lut[1597] = 662;  
        func_lut[1598] = 660;  
        func_lut[1599] = 658;  
        func_lut[1600] = 657;  
        func_lut[1601] = 655;  
        func_lut[1602] = 653;  
        func_lut[1603] = 652;  
        func_lut[1604] = 650;  
        func_lut[1605] = 649;  
        func_lut[1606] = 647;  
        func_lut[1607] = 645;  
        func_lut[1608] = 644;  
        func_lut[1609] = 642;  
        func_lut[1610] = 641;  
        func_lut[1611] = 639;  
        func_lut[1612] = 637;  
        func_lut[1613] = 636;  
        func_lut[1614] = 634;  
        func_lut[1615] = 633;  
        func_lut[1616] = 631;  
        func_lut[1617] = 630;  
        func_lut[1618] = 628;  
        func_lut[1619] = 627;  
        func_lut[1620] = 625;  
        func_lut[1621] = 624;  
        func_lut[1622] = 622;  
        func_lut[1623] = 621;  
        func_lut[1624] = 619;  
        func_lut[1625] = 618;  
        func_lut[1626] = 616;  
        func_lut[1627] = 615;  
        func_lut[1628] = 613;  
        func_lut[1629] = 612;  
        func_lut[1630] = 610;  
        func_lut[1631] = 609;  
        func_lut[1632] = 607;  
        func_lut[1633] = 606;  
        func_lut[1634] = 604;  
        func_lut[1635] = 603;  
        func_lut[1636] = 602;  
        func_lut[1637] = 600;  
        func_lut[1638] = 599;  
        func_lut[1639] = 597;  
        func_lut[1640] = 596;  
        func_lut[1641] = 594;  
        func_lut[1642] = 593;  
        func_lut[1643] = 592;  
        func_lut[1644] = 590;  
        func_lut[1645] = 589;  
        func_lut[1646] = 587;  
        func_lut[1647] = 586;  
        func_lut[1648] = 585;  
        func_lut[1649] = 583;  
        func_lut[1650] = 582;  
        func_lut[1651] = 581;  
        func_lut[1652] = 579;  
        func_lut[1653] = 578;  
        func_lut[1654] = 577;  
        func_lut[1655] = 575;  
        func_lut[1656] = 574;  
        func_lut[1657] = 573;  
        func_lut[1658] = 571;  
        func_lut[1659] = 570;  
        func_lut[1660] = 569;  
        func_lut[1661] = 567;  
        func_lut[1662] = 566;  
        func_lut[1663] = 565;  
        func_lut[1664] = 563;  
        func_lut[1665] = 562;  
        func_lut[1666] = 561;  
        func_lut[1667] = 559;  
        func_lut[1668] = 558;  
        func_lut[1669] = 557;  
        func_lut[1670] = 556;  
        func_lut[1671] = 554;  
        func_lut[1672] = 553;  
        func_lut[1673] = 552;  
        func_lut[1674] = 551;  
        func_lut[1675] = 549;  
        func_lut[1676] = 548;  
        func_lut[1677] = 547;  
        func_lut[1678] = 546;  
        func_lut[1679] = 544;  
        func_lut[1680] = 543;  
        func_lut[1681] = 542;  
        func_lut[1682] = 541;  
        func_lut[1683] = 539;  
        func_lut[1684] = 538;  
        func_lut[1685] = 537;  
        func_lut[1686] = 536;  
        func_lut[1687] = 535;  
        func_lut[1688] = 533;  
        func_lut[1689] = 532;  
        func_lut[1690] = 531;  
        func_lut[1691] = 530;  
        func_lut[1692] = 529;  
        func_lut[1693] = 528;  
        func_lut[1694] = 526;  
        func_lut[1695] = 525;  
        func_lut[1696] = 524;  
        func_lut[1697] = 523;  
        func_lut[1698] = 522;  
        func_lut[1699] = 521;  
        func_lut[1700] = 519;  
        func_lut[1701] = 518;  
        func_lut[1702] = 517;  
        func_lut[1703] = 516;  
        func_lut[1704] = 515;  
        func_lut[1705] = 514;  
        func_lut[1706] = 513;  
        func_lut[1707] = 511;  
        func_lut[1708] = 510;  
        func_lut[1709] = 509;  
        func_lut[1710] = 508;  
        func_lut[1711] = 507;  
        func_lut[1712] = 506;  
        func_lut[1713] = 505;  
        func_lut[1714] = 504;  
        func_lut[1715] = 503;  
        func_lut[1716] = 501;  
        func_lut[1717] = 500;  
        func_lut[1718] = 499;  
        func_lut[1719] = 498;  
        func_lut[1720] = 497;  
        func_lut[1721] = 496;  
        func_lut[1722] = 495;  
        func_lut[1723] = 494;  
        func_lut[1724] = 493;  
        func_lut[1725] = 492;  
        func_lut[1726] = 491;  
        func_lut[1727] = 490;  
        func_lut[1728] = 489;  
        func_lut[1729] = 488;  
        func_lut[1730] = 487;  
        func_lut[1731] = 485;  
        func_lut[1732] = 484;  
        func_lut[1733] = 483;  
        func_lut[1734] = 482;  
        func_lut[1735] = 481;  
        func_lut[1736] = 480;  
        func_lut[1737] = 479;  
        func_lut[1738] = 478;  
        func_lut[1739] = 477;  
        func_lut[1740] = 476;  
        func_lut[1741] = 475;  
        func_lut[1742] = 474;  
        func_lut[1743] = 473;  
        func_lut[1744] = 472;  
        func_lut[1745] = 471;  
        func_lut[1746] = 470;  
        func_lut[1747] = 469;  
        func_lut[1748] = 468;  
        func_lut[1749] = 467;  
        func_lut[1750] = 466;  
        func_lut[1751] = 465;  
        func_lut[1752] = 464;  
        func_lut[1753] = 463;  
        func_lut[1754] = 462;  
        func_lut[1755] = 461;  
        func_lut[1756] = 461;  
        func_lut[1757] = 460;  
        func_lut[1758] = 459;  
        func_lut[1759] = 458;  
        func_lut[1760] = 457;  
        func_lut[1761] = 456;  
        func_lut[1762] = 455;  
        func_lut[1763] = 454;  
        func_lut[1764] = 453;  
        func_lut[1765] = 452;  
        func_lut[1766] = 451;  
        func_lut[1767] = 450;  
        func_lut[1768] = 449;  
        func_lut[1769] = 448;  
        func_lut[1770] = 447;  
        func_lut[1771] = 446;  
        func_lut[1772] = 446;  
        func_lut[1773] = 445;  
        func_lut[1774] = 444;  
        func_lut[1775] = 443;  
        func_lut[1776] = 442;  
        func_lut[1777] = 441;  
        func_lut[1778] = 440;  
        func_lut[1779] = 439;  
        func_lut[1780] = 438;  
        func_lut[1781] = 437;  
        func_lut[1782] = 437;  
        func_lut[1783] = 436;  
        func_lut[1784] = 435;  
        func_lut[1785] = 434;  
        func_lut[1786] = 433;  
        func_lut[1787] = 432;  
        func_lut[1788] = 431;  
        func_lut[1789] = 430;  
        func_lut[1790] = 430;  
        func_lut[1791] = 429;  
        func_lut[1792] = 428;  
        func_lut[1793] = 427;  
        func_lut[1794] = 426;  
        func_lut[1795] = 425;  
        func_lut[1796] = 424;  
        func_lut[1797] = 424;  
        func_lut[1798] = 423;  
        func_lut[1799] = 422;  
        func_lut[1800] = 421;  
        func_lut[1801] = 420;  
        func_lut[1802] = 419;  
        func_lut[1803] = 419;  
        func_lut[1804] = 418;  
        func_lut[1805] = 417;  
        func_lut[1806] = 416;  
        func_lut[1807] = 415;  
        func_lut[1808] = 414;  
        func_lut[1809] = 414;  
        func_lut[1810] = 413;  
        func_lut[1811] = 412;  
        func_lut[1812] = 411;  
        func_lut[1813] = 410;  
        func_lut[1814] = 410;  
        func_lut[1815] = 409;  
        func_lut[1816] = 408;  
        func_lut[1817] = 407;  
        func_lut[1818] = 406;  
        func_lut[1819] = 406;  
        func_lut[1820] = 405;  
        func_lut[1821] = 404;  
        func_lut[1822] = 403;  
        func_lut[1823] = 402;  
        func_lut[1824] = 402;  
        func_lut[1825] = 401;  
        func_lut[1826] = 400;  
        func_lut[1827] = 399;  
        func_lut[1828] = 398;  
        func_lut[1829] = 398;  
        func_lut[1830] = 397;  
        func_lut[1831] = 396;  
        func_lut[1832] = 395;  
        func_lut[1833] = 395;  
        func_lut[1834] = 394;  
        func_lut[1835] = 393;  
        func_lut[1836] = 392;  
        func_lut[1837] = 392;  
        func_lut[1838] = 391;  
        func_lut[1839] = 390;  
        func_lut[1840] = 389;  
        func_lut[1841] = 389;  
        func_lut[1842] = 388;  
        func_lut[1843] = 387;  
        func_lut[1844] = 386;  
        func_lut[1845] = 386;  
        func_lut[1846] = 385;  
        func_lut[1847] = 384;  
        func_lut[1848] = 383;  
        func_lut[1849] = 383;  
        func_lut[1850] = 382;  
        func_lut[1851] = 381;  
        func_lut[1852] = 381;  
        func_lut[1853] = 380;  
        func_lut[1854] = 379;  
        func_lut[1855] = 378;  
        func_lut[1856] = 378;  
        func_lut[1857] = 377;  
        func_lut[1858] = 376;  
        func_lut[1859] = 376;  
        func_lut[1860] = 375;  
        func_lut[1861] = 374;  
        func_lut[1862] = 373;  
        func_lut[1863] = 373;  
        func_lut[1864] = 372;  
        func_lut[1865] = 371;  
        func_lut[1866] = 371;  
        func_lut[1867] = 370;  
        func_lut[1868] = 369;  
        func_lut[1869] = 369;  
        func_lut[1870] = 368;  
        func_lut[1871] = 367;  
        func_lut[1872] = 367;  
        func_lut[1873] = 366;  
        func_lut[1874] = 365;  
        func_lut[1875] = 365;  
        func_lut[1876] = 364;  
        func_lut[1877] = 363;  
        func_lut[1878] = 363;  
        func_lut[1879] = 362;  
        func_lut[1880] = 361;  
        func_lut[1881] = 361;  
        func_lut[1882] = 360;  
        func_lut[1883] = 359;  
        func_lut[1884] = 359;  
        func_lut[1885] = 358;  
        func_lut[1886] = 357;  
        func_lut[1887] = 357;  
        func_lut[1888] = 356;  
        func_lut[1889] = 355;  
        func_lut[1890] = 355;  
        func_lut[1891] = 354;  
        func_lut[1892] = 353;  
        func_lut[1893] = 353;  
        func_lut[1894] = 352;  
        func_lut[1895] = 351;  
        func_lut[1896] = 351;  
        func_lut[1897] = 350;  
        func_lut[1898] = 349;  
        func_lut[1899] = 349;  
        func_lut[1900] = 348;  
        func_lut[1901] = 348;  
        func_lut[1902] = 347;  
        func_lut[1903] = 346;  
        func_lut[1904] = 346;  
        func_lut[1905] = 345;  
        func_lut[1906] = 344;  
        func_lut[1907] = 344;  
        func_lut[1908] = 343;  
        func_lut[1909] = 343;  
        func_lut[1910] = 342;  
        func_lut[1911] = 341;  
        func_lut[1912] = 341;  
        func_lut[1913] = 340;  
        func_lut[1914] = 340;  
        func_lut[1915] = 339;  
        func_lut[1916] = 338;  
        func_lut[1917] = 338;  
        func_lut[1918] = 337;  
        func_lut[1919] = 337;  
        func_lut[1920] = 336;  
        func_lut[1921] = 335;  
        func_lut[1922] = 335;  
        func_lut[1923] = 334;  
        func_lut[1924] = 334;  
        func_lut[1925] = 333;  
        func_lut[1926] = 332;  
        func_lut[1927] = 332;  
        func_lut[1928] = 331;  
        func_lut[1929] = 331;  
        func_lut[1930] = 330;  
        func_lut[1931] = 329;  
        func_lut[1932] = 329;  
        func_lut[1933] = 328;  
        func_lut[1934] = 328;  
        func_lut[1935] = 327;  
        func_lut[1936] = 327;  
        func_lut[1937] = 326;  
        func_lut[1938] = 325;  
        func_lut[1939] = 325;  
        func_lut[1940] = 324;  
        func_lut[1941] = 324;  
        func_lut[1942] = 323;  
        func_lut[1943] = 323;  
        func_lut[1944] = 322;  
        func_lut[1945] = 321;  
        func_lut[1946] = 321;  
        func_lut[1947] = 320;  
        func_lut[1948] = 320;  
        func_lut[1949] = 319;  
        func_lut[1950] = 319;  
        func_lut[1951] = 318;  
        func_lut[1952] = 318;  
        func_lut[1953] = 317;  
        func_lut[1954] = 316;  
        func_lut[1955] = 316;  
        func_lut[1956] = 315;  
        func_lut[1957] = 315;  
        func_lut[1958] = 314;  
        func_lut[1959] = 314;  
        func_lut[1960] = 313;  
        func_lut[1961] = 313;  
        func_lut[1962] = 312;  
        func_lut[1963] = 312;  
        func_lut[1964] = 311;  
        func_lut[1965] = 311;  
        func_lut[1966] = 310;  
        func_lut[1967] = 309;  
        func_lut[1968] = 309;  
        func_lut[1969] = 308;  
        func_lut[1970] = 308;  
        func_lut[1971] = 307;  
        func_lut[1972] = 307;  
        func_lut[1973] = 306;  
        func_lut[1974] = 306;  
        func_lut[1975] = 305;  
        func_lut[1976] = 305;  
        func_lut[1977] = 304;  
        func_lut[1978] = 304;  
        func_lut[1979] = 303;  
        func_lut[1980] = 303;  
        func_lut[1981] = 302;  
        func_lut[1982] = 302;  
        func_lut[1983] = 301;  
        func_lut[1984] = 301;  
        func_lut[1985] = 300;  
        func_lut[1986] = 300;  
        func_lut[1987] = 299;  
        func_lut[1988] = 299;  
        func_lut[1989] = 298;  
        func_lut[1990] = 298;  
        func_lut[1991] = 297;  
        func_lut[1992] = 297;  
        func_lut[1993] = 296;  
        func_lut[1994] = 296;  
        func_lut[1995] = 295;  
        func_lut[1996] = 295;  
        func_lut[1997] = 294;  
        func_lut[1998] = 294;  
        func_lut[1999] = 293;  
        func_lut[2000] = 293;  
        func_lut[2001] = 292;  
        func_lut[2002] = 292;  
        func_lut[2003] = 291;  
        func_lut[2004] = 291;  
        func_lut[2005] = 290;  
        func_lut[2006] = 290;  
        func_lut[2007] = 289;  
        func_lut[2008] = 289;  
        func_lut[2009] = 288;  
        func_lut[2010] = 288;  
        func_lut[2011] = 287;  
        func_lut[2012] = 287;  
        func_lut[2013] = 287;  
        func_lut[2014] = 286;  
        func_lut[2015] = 286;  
        func_lut[2016] = 285;  
        func_lut[2017] = 285;  
        func_lut[2018] = 284;  
        func_lut[2019] = 284;  
        func_lut[2020] = 283;  
        func_lut[2021] = 283;  
        func_lut[2022] = 282;  
        func_lut[2023] = 282;  
        func_lut[2024] = 281;  
        func_lut[2025] = 281;  
        func_lut[2026] = 281;  
        func_lut[2027] = 280;  
        func_lut[2028] = 280;  
        func_lut[2029] = 279;  
        func_lut[2030] = 279;  
        func_lut[2031] = 278;  
        func_lut[2032] = 278;  
        func_lut[2033] = 277;  
        func_lut[2034] = 277;  
        func_lut[2035] = 276;  
        func_lut[2036] = 276;  
        func_lut[2037] = 276;  
        func_lut[2038] = 275;  
        func_lut[2039] = 275;  
        func_lut[2040] = 274;  
        func_lut[2041] = 274;  
        func_lut[2042] = 273;  
        func_lut[2043] = 273;  
        func_lut[2044] = 272;  
        func_lut[2045] = 272;  
        func_lut[2046] = 272;  
        func_lut[2047] = 271; 
    end

endmodule